* /home/fossee/Downloads/powercktexamples/fullwaverec/fullwaverec.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Dec  4 15:43:40 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
x1  GND pulse out2 SCR		
v1  in1 in2 sine		
v2  pulse GND pulse		
D1  in1 out1 D		
D3  in2 out1 D		
D2  GND in1 D		
D4  GND in2 D		
R1  out1 out2 100		

.end
