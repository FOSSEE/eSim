* C:\FOSSEE\eSim\library\SubcircuitLibrary\14_lm386\14_lm386.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/14/25 17:23:21

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q2  Net-_Q2-Pad1_ Net-_Q1-Pad3_ Net-_Q2-Pad3_ eSim_PNP		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_PNP		
Q3  Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_Q1-Pad1_ eSim_NPN		
Q5  Net-_Q4-Pad1_ Net-_Q5-Pad2_ Net-_Q5-Pad3_ eSim_PNP		
Q4  Net-_Q4-Pad1_ Net-_Q2-Pad1_ Net-_Q1-Pad1_ eSim_NPN		
Q6  Net-_Q1-Pad1_ Net-_Q6-Pad2_ Net-_Q5-Pad2_ eSim_PNP		
Q7  Net-_D2-Pad2_ Net-_Q4-Pad1_ Net-_Q1-Pad1_ eSim_NPN		
Q8  Net-_Q10-Pad2_ Net-_D2-Pad2_ Net-_Q10-Pad1_ eSim_PNP		
Q10  Net-_Q10-Pad1_ Net-_Q10-Pad2_ Net-_Q1-Pad1_ eSim_NPN		
R1  Net-_Q1-Pad2_ Net-_Q1-Pad1_ 50k		
R4  Net-_Q2-Pad3_ Net-_R4-Pad2_ 150		
R5  Net-_R4-Pad2_ Net-_Q5-Pad3_ 1.35k		
R6  Net-_Q5-Pad3_ Net-_Q10-Pad1_ 15k		
R3  Net-_R2-Pad2_ Net-_Q2-Pad3_ 15k		
R2  Net-_Q9-Pad1_ Net-_R2-Pad2_ 15k		
R7  Net-_Q6-Pad2_ Net-_Q1-Pad1_ 50k		
D2  Net-_D1-Pad2_ Net-_D2-Pad2_ eSim_Diode		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
R8  Net-_Q9-Pad1_ Net-_D1-Pad1_ 1.35k		
Q9  Net-_Q9-Pad1_ Net-_D1-Pad1_ Net-_Q10-Pad1_ eSim_NPN		
U1  Net-_Q5-Pad3_ Net-_Q1-Pad2_ Net-_Q6-Pad2_ Net-_Q1-Pad1_ Net-_Q10-Pad1_ Net-_Q9-Pad1_ Net-_R2-Pad2_ Net-_R4-Pad2_ PORT		

.end
