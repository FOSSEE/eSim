* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Jun  8 12:02:52 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
v1  6 0 DC		
v2  2 0 AC		
R1  3 2 50		
R2  6 8 200k		
C1  3 8 40u		
R3  8 0 50k		
R6  4 0 1k		
C2  0 5 100u		
C3  4 7 40u		
R5  6 7 2k		
R4  5 0 1.5k		
Q1  7 8 5 NPN		

.end
