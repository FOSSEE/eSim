.title KiCad schematic
Q6 Net-_Q1-Pad3_ Net-_Q6-Pad2_ Net-_Q5-Pad3_ eSim_NPN
R4 Net-_Q1-Pad3_ Net-_C1-Pad1_ 200k
U3 Net-_Q5-Pad2_ Net-_Q6-Pad2_ GND Net-_Q12-Pad3_ Net-_Q12-Pad3_ Net-_Q10-Pad3_ Net-_Q6-Pad2_ Net-_Q5-Pad2_ PORT
R6 GND Net-_Q7-Pad3_ 47k
Q7 Net-_Q7-Pad1_ Net-_C1-Pad1_ Net-_Q7-Pad3_ eSim_NPN
Q13 Net-_Q10-Pad3_ Net-_C1-Pad2_ Net-_Q13-Pad3_ eSim_NPN
Q10 Net-_C1-Pad2_ Net-_Q10-Pad2_ Net-_Q10-Pad3_ eSim_PNP
R8 Net-_Q12-Pad2_ Net-_Q13-Pad3_ 4.7k
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ eSim_Diode
D3 Net-_D2-Pad2_ GND eSim_Diode
R5 GND Net-_Q5-Pad3_ 10k
Q5 Net-_C1-Pad1_ Net-_Q5-Pad2_ Net-_Q5-Pad3_ eSim_NPN
U1 GND Net-_D1-Pad1_ zener
Q2 GND Net-_Q1-Pad1_ Net-_Q10-Pad2_ eSim_PNP
R1 Net-_D1-Pad1_ Net-_Q10-Pad3_ 250k
U2 GND Net-_D1-Pad2_ zener
R3 Net-_Q5-Pad2_ Net-_D2-Pad1_ 250k
R2 Net-_D2-Pad1_ Net-_Q1-Pad3_ 100k
Q1 Net-_Q1-Pad1_ Net-_D1-Pad2_ Net-_Q1-Pad3_ eSim_NPN
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode
R7 GND Net-_Q11-Pad2_ 47k
Q9 Net-_Q7-Pad1_ Net-_Q7-Pad3_ Net-_Q11-Pad2_ eSim_NPN
Q11 Net-_C1-Pad2_ Net-_Q11-Pad2_ GND eSim_NPN
Q12 Net-_C1-Pad2_ Net-_Q12-Pad2_ Net-_Q12-Pad3_ eSim_NPN
Q15 Net-_Q12-Pad3_ Net-_Q11-Pad2_ GND eSim_NPN
R9 Net-_Q12-Pad3_ Net-_Q12-Pad2_ 50k
Q14 Net-_Q10-Pad3_ Net-_Q13-Pad3_ Net-_Q12-Pad2_ eSim_NPN
Q3 Net-_Q1-Pad1_ Net-_Q3-Pad2_ Net-_Q10-Pad3_ eSim_PNP
Q4 Net-_D1-Pad2_ Net-_Q1-Pad1_ Net-_Q3-Pad2_ eSim_PNP
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 1uf
Q8 Net-_Q10-Pad3_ Net-_D1-Pad2_ Net-_Q7-Pad1_ eSim_NPN
.end
