.title KiCad schematic
v1 Net-_M2-Pad1_ GND 5
U10 Net-_M1-Pad1_ Net-_U1-Pad3_ adc_bridge_1
U1 Net-_U1-Pad1_ Net-_U3-Pad1_ Net-_U1-Pad3_ PORT
U9 Net-_U7-Pad3_ Net-_M2-Pad2_ dac_bridge_1
U11 Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ d_and
M2 Net-_M2-Pad1_ Net-_M2-Pad2_ Net-_M1-Pad1_ Net-_M2-Pad1_ eSim_MOS_P
M1 Net-_M1-Pad1_ Net-_M1-Pad2_ GND GND eSim_MOS_N
U12 Net-_U11-Pad3_ Net-_M1-Pad2_ dac_bridge_1
U6 Net-_U4-Pad2_ Net-_U11-Pad1_ d_inverter
U7 Net-_U3-Pad2_ Net-_U4-Pad2_ Net-_U7-Pad3_ d_nand
U8 Net-_U5-Pad2_ Net-_U11-Pad2_ d_inverter
U5 Net-_U3-Pad2_ Net-_U5-Pad2_ d_inverter
U4 Net-_U2-Pad2_ Net-_U4-Pad2_ d_inverter
U3 Net-_U3-Pad1_ Net-_U3-Pad2_ d_inverter
U2 Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter
.end
