* E:\IC_811M\IC_811M.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/09/25 21:52:29

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R2-Pad2_ Net-_R1-Pad2_ Net-_X1-Pad3_ GND ? OUT Net-_X1-Pad7_ GND GND GND TL811M		
R1  IN Net-_R1-Pad2_ 50k		
R2  IN Net-_R2-Pad2_ 50k		
v2  Net-_X1-Pad7_ GND DC		
v3  Net-_X1-Pad3_ GND DC		
U1  OUT plot_v1		
U2  IN plot_v1		
v1  IN GND pulse		

.end
