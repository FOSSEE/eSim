* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Jun 12 12:25:06 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
C1  3 4 1u		
v1  1 4 dc		
v2  2 4 5		
M1  3 1 4 4 MOS_N		
M2  3 1 2 2 MOS_P		

.end
