* C:\FOSSEE\eSim\library\SubcircuitLibrary\74HC20\74HC20.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/13/25 16:05:56

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U10-Pad1_ d_inverter		
U3  Net-_U1-Pad2_ Net-_U10-Pad2_ d_inverter		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ d_nor		
U4  Net-_U1-Pad3_ Net-_U11-Pad1_ d_inverter		
U5  Net-_U1-Pad4_ Net-_U11-Pad2_ d_inverter		
U11  Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ d_nor		
U14  Net-_U10-Pad3_ Net-_U11-Pad3_ Net-_U14-Pad3_ d_nand		
U16  Net-_U14-Pad3_ Net-_U16-Pad2_ d_inverter		
U18  Net-_U16-Pad2_ Net-_U1-Pad5_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ PORT		
U6  Net-_U1-Pad6_ Net-_U12-Pad1_ d_inverter		
U7  Net-_U1-Pad7_ Net-_U12-Pad2_ d_inverter		
U12  Net-_U12-Pad1_ Net-_U12-Pad2_ Net-_U12-Pad3_ d_nor		
U8  Net-_U1-Pad8_ Net-_U13-Pad1_ d_inverter		
U9  Net-_U1-Pad9_ Net-_U13-Pad2_ d_inverter		
U13  Net-_U13-Pad1_ Net-_U13-Pad2_ Net-_U13-Pad3_ d_nor		
U15  Net-_U12-Pad3_ Net-_U13-Pad3_ Net-_U15-Pad3_ d_nand		
U17  Net-_U15-Pad3_ Net-_U17-Pad2_ d_inverter		
U19  Net-_U17-Pad2_ Net-_U1-Pad10_ d_inverter		

.end
