.title KiCad schematic
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ eSim_Diode
Q6 Net-_Q4-Pad1_ Net-_D2-Pad2_ Net-_D3-Pad2_ eSim_PNP
Q7 Net-_D4-Pad1_ Net-_D6-Pad2_ Net-_D3-Pad1_ eSim_PNP
Q2 Net-_D2-Pad1_ Net-_D3-Pad2_ Net-_D3-Pad1_ eSim_PNP
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ eSim_Diode
Q4 Net-_Q4-Pad1_ Net-_D2-Pad1_ Net-_D2-Pad2_ eSim_PNP
U1 Net-_Q10-Pad1_ Net-_Q1-Pad2_ Net-_Q5-Pad2_ Net-_D1-Pad2_ Net-_D1-Pad1_ Net-_Q13-Pad3_ Net-_D3-Pad1_ Net-_Q13-Pad1_ PORT
Q5 Net-_D4-Pad1_ Net-_Q5-Pad2_ Net-_Q1-Pad3_ eSim_NPN
Q1 Net-_D2-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode
Q3 Net-_Q1-Pad3_ Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_NPN
Q8 Net-_Q4-Pad1_ Net-_D5-Pad1_ Net-_D1-Pad2_ eSim_NPN
Q12 Net-_Q12-Pad1_ Net-_Q10-Pad1_ Net-_Q12-Pad3_ eSim_NPN
Q9 Net-_Q10-Pad1_ Net-_Q4-Pad1_ Net-_D5-Pad1_ eSim_NPN
D5 Net-_D5-Pad1_ Net-_D1-Pad2_ eSim_Diode
R2 Net-_Q13-Pad3_ Net-_Q12-Pad3_ 47k
Q13 Net-_Q13-Pad1_ Net-_Q12-Pad3_ Net-_Q13-Pad3_ eSim_NPN
D4 Net-_D4-Pad1_ Net-_D4-Pad2_ eSim_Diode
R1 Net-_Q12-Pad1_ Net-_D3-Pad1_ 2k
D6 Net-_D3-Pad1_ Net-_D6-Pad2_ eSim_Diode
Q10 Net-_Q10-Pad1_ Net-_D4-Pad1_ Net-_D4-Pad2_ eSim_PNP
Q11 Net-_Q10-Pad1_ Net-_D4-Pad2_ Net-_D6-Pad2_ eSim_PNP
.end
