* C:\FOSSEE\eSim\library\SubcircuitLibrary\XOR\XOR.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/28/24 11:19:17

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M1-Pad3_ Net-_M2-Pad2_ GND GND mosfet_n		
M8  Net-_M7-Pad3_ Net-_M6-Pad2_ GND GND mosfet_n		
M7  Net-_M1-Pad1_ Net-_M4-Pad2_ Net-_M7-Pad3_ Net-_M7-Pad3_ mosfet_n		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_n		
M4  Net-_M3-Pad3_ Net-_M4-Pad2_ Net-_M1-Pad1_ Net-_M3-Pad3_ mosfet_p		
M6  Net-_M3-Pad3_ Net-_M6-Pad2_ Net-_M1-Pad1_ Net-_M3-Pad3_ mosfet_p		
M3  Net-_M3-Pad1_ Net-_M1-Pad2_ Net-_M3-Pad3_ Net-_M3-Pad1_ mosfet_p		
M5  Net-_M3-Pad1_ Net-_M2-Pad2_ Net-_M3-Pad3_ Net-_M3-Pad1_ mosfet_p		
X1  Net-_M1-Pad2_ Net-_M4-Pad2_ NOT_Gate		
X2  Net-_M2-Pad2_ Net-_M6-Pad2_ NOT_Gate		
v1  Net-_M3-Pad1_ GND DC		
U1  Net-_M1-Pad2_ Net-_M2-Pad2_ Net-_M1-Pad1_ PORT		

.end
