* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/TFF_SR/TFF_SR.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jul  9 11:21:42 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad2_ Net-_U1-Pad8_ Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_X1-Pad5_ Net-_U1-Pad3_ NAND_3		
X3  Net-_U1-Pad5_ Net-_X1-Pad5_ Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad7_ Net-_U1-Pad8_ NAND_3		
X2  Net-_U1-Pad3_ Net-_U1-Pad7_ Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_X2-Pad5_ Net-_U1-Pad2_ NAND_3		
X4  Net-_U1-Pad7_ Net-_X2-Pad5_ Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad8_ Net-_U1-Pad6_ NAND_3		
scmode1  SKY130mode		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ PORT		

.end
