.title KiCad schematic
U3 K plot_v1
U2 CLK plot_v1
U1 J plot_v1
Vk1 K GND DC
Vj1 J GND DC
Vclk1 CLK GND pulse
Vclr1 Net-_U4-Pad3_ GND DC
Vcc1 Net-_Vcc1-Pad1_ GND 5
X1 Net-_U4-Pad6_ Net-_U4-Pad7_ Net-_U4-Pad8_ Net-_Vcc1-Pad1_ unconnected-_X1-Pad5_ unconnected-_X1-Pad6_ unconnected-_X1-Pad7_ unconnected-_X1-Pad8_ unconnected-_X1-Pad9_ unconnected-_X1-Pad10_ GND Net-_U7-Pad1_ Net-_U7-Pad2_ Net-_U4-Pad5_ SN5473
U6 NQ plot_v1
U4 J CLK Net-_U4-Pad3_ K Net-_U4-Pad5_ Net-_U4-Pad6_ Net-_U4-Pad7_ Net-_U4-Pad8_ adc_bridge_4
U5 Q plot_v1
U7 Net-_U7-Pad1_ Net-_U7-Pad2_ Q NQ dac_bridge_2
R2 GND NQ 1k
R1 GND Q 1k
.end
