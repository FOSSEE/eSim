* C:\FOSSEE\eSim\library\SubcircuitLibrary\NAND\NAND.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/25/24 01:53:20

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M2-Pad3_ Net-_M3-Pad2_ GND GND mosfet_n		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M4  Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M2  Net-_M1-Pad3_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_n		
v1  Net-_M1-Pad1_ GND DC		
U1  Net-_M1-Pad2_ Net-_M3-Pad2_ Net-_M1-Pad3_ PORT		

.end
