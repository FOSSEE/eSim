* C:\FOSSEE\eSim\library\SubcircuitLibrary\mux4\mux4.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/02/25 13:58:33

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter		
U3  Net-_U1-Pad2_ Net-_U3-Pad2_ d_inverter		
X1  Net-_U2-Pad2_ Net-_U3-Pad2_ Net-_U1-Pad6_ Net-_X1-Pad4_ 3_and		
X2  Net-_U1-Pad1_ Net-_U3-Pad2_ Net-_U1-Pad3_ Net-_X2-Pad4_ 3_and		
X3  Net-_U2-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad4_ Net-_X3-Pad4_ 3_and		
X4  Net-_U1-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad5_ Net-_X4-Pad4_ 3_and		
X5  Net-_X1-Pad4_ Net-_X2-Pad4_ Net-_X3-Pad4_ Net-_X4-Pad4_ Net-_U1-Pad7_ 4_OR		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ PORT		

.end
