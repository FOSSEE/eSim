* C:\FOSSEE\eSim\library\SubcircuitLibrary\CD4027B_IC\CD4027B_IC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/29/24 12:20:01

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad15_ Net-_U1-Pad14_ Net-_U1-Pad16_ Net-_U1-Pad8_ JK_FF		
X2  Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad5_ Net-_U1-Pad4_ Net-_U1-Pad3_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad16_ Net-_U1-Pad8_ JK_FF		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ PORT		

.end
