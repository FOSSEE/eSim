.title KiCad schematic
U6 Net-_V_OEn1-Pad1_ Net-_V_A0-Pad1_ Net-_V_A1-Pad1_ Net-_V_A2-Pad1_ Net-_V_A3-Pad1_ Net-_U6-Pad6_ Net-_U6-Pad7_ Net-_U6-Pad8_ Net-_U6-Pad9_ Net-_U6-Pad10_ adc_bridge_5
V_OEn1 Net-_V_OEn1-Pad1_ GND DC
V_A3 Net-_V_A3-Pad1_ GND DC
U5 Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ V_A4 V_A5 V_A6 V_A7 dac_bridge_4
U1 V_A4 plot_v1
U3 V_A6 plot_v1
U4 V_A7 plot_v1
U2 V_A5 plot_v1
v1 Net-_v1-Pad1_ GND 5
U7 Net-_V_DIR1-Pad1_ Net-_U7-Pad2_ adc_bridge_1
U8 Net-_U8-Pad1_ Net-_U8-Pad2_ Net-_U8-Pad3_ Net-_U8-Pad4_ V_B0 V_B1 V_B2 V_B3 dac_bridge_4
U9 Net-_V_B4-Pad1_ Net-_V_5-Pad1_ Net-_V_B6-Pad1_ Net-_V_B7-Pad1_ Net-_U9-Pad5_ Net-_U9-Pad6_ Net-_U9-Pad7_ Net-_U9-Pad8_ adc_bridge_4
X1 Net-_U6-Pad6_ Net-_U6-Pad7_ Net-_U6-Pad8_ Net-_U6-Pad9_ Net-_U6-Pad10_ Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U5-Pad3_ Net-_U5-Pad4_ GND Net-_U9-Pad8_ Net-_U9-Pad7_ Net-_U9-Pad6_ Net-_U9-Pad5_ Net-_U8-Pad4_ Net-_U8-Pad3_ Net-_U8-Pad2_ Net-_U8-Pad1_ Net-_U7-Pad2_ Net-_v1-Pad1_ 74HC245
V_B7 Net-_V_B7-Pad1_ GND DC
V_B6 Net-_V_B6-Pad1_ GND DC
V_DIR1 Net-_V_DIR1-Pad1_ GND DC
U11 V_B1 plot_v1
U12 V_B2 plot_v1
U13 V_B3 plot_v1
U10 V_B0 plot_v1
V_5 Net-_V_5-Pad1_ GND DC
V_B4 Net-_V_B4-Pad1_ GND DC
V_A0 Net-_V_A0-Pad1_ GND DC
V_A2 Net-_V_A2-Pad1_ GND DC
V_A1 Net-_V_A1-Pad1_ GND DC
.end
