* /home/bhargav/Downloads/eSim-1.1.2/src/SubcircuitLibrary/IB3858/IB3858.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Jun 24 16:30:15 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  Net-_R1-Pad1_ Net-_L1-Pad1_ 5.2		
L1  Net-_L1-Pad1_ Net-_C1-Pad1_ 3.08m		
L2  Net-_C1-Pad1_ Net-_C1-Pad2_ 61.100458m		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 896.8481u		
R2  Net-_C1-Pad1_ Net-_C1-Pad2_ 73.6254		
U1  Net-_R1-Pad1_ Net-_C1-Pad2_ PORT		

.end
