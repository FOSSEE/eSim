* C:\Users\Shanthipriya\eSim-Workspace\030\030.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/29/25 13:20:44

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U9-Pad9_ Net-_U9-Pad10_ Net-_U9-Pad11_ Net-_U9-Pad12_ Net-_U9-Pad13_ Net-_U9-Pad14_ Net-_U9-Pad15_ Net-_U9-Pad16_ Net-_U10-Pad1_ 74_1030		
U9  A1 A2 A3 A4 A5 A6 A7 A8 Net-_U9-Pad9_ Net-_U9-Pad10_ Net-_U9-Pad11_ Net-_U9-Pad12_ Net-_U9-Pad13_ Net-_U9-Pad14_ Net-_U9-Pad15_ Net-_U9-Pad16_ adc_bridge_8		
U10  Net-_U10-Pad1_ OUT dac_bridge_1		
v1  A1 GND pulse		
v2  A2 GND pulse		
v3  A3 GND pulse		
v4  A4 GND pulse		
v5  A5 GND pulse		
v6  A6 GND pulse		
v7  A7 GND pulse		
v8  A8 GND pulse		
U11  OUT plot_v1		
U1  A1 plot_v1		
U2  A2 plot_v1		
U3  A3 plot_v1		
U4  A4 plot_v1		
U5  A5 plot_v1		
U6  A6 plot_v1		
U7  A7 plot_v1		
U8  A8 plot_v1		

.end
