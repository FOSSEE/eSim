* C:\Users\Aditya\eSim-Workspace\9348\9348.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/03/24 16:25:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v2  Net-_X1-Pad16_ GND DC		
R1  PO GND 1000k		
R2  PE GND 1000k		
X1  i5 i6 i7 i8 i9 i10 i11 GND PO PE i0 i1 i2 i3 i4 Net-_X1-Pad16_ 9348_IC		
U2  PE plot_v1		
U1  PO plot_v1		
v1  i5 GND pulse		
v3  i6 GND pulse		
v4  i7 GND pulse		
v5  i8 GND pulse		
v6  i9 GND pulse		
v7  i10 GND pulse		
v8  i11 GND pulse		
v9  i0 GND pulse		
v10  i1 GND pulse		
v11  i2 GND pulse		
v12  i3 GND pulse		
v13  i4 GND pulse		
U4  i6 plot_v1		
U5  i7 plot_v1		
U6  i8 plot_v1		
U7  i9 plot_v1		
U8  i10 plot_v1		
U9  i11 plot_v1		
U10  i0 plot_v1		
U11  i1 plot_v1		
U12  i2 plot_v1		
U13  i3 plot_v1		
U14  i4 plot_v1		
U3  i5 plot_v1		

.end
