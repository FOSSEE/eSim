* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 26 October 2015 03:08:36 PM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
v1  1 0 DC		
R1  1 2 1k		
D1  2 0 D		

.end
