* C:\FOSSEE\eSim\library\SubcircuitLibrary\74688\74688.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/21/25 17:00:02

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter		
U3  Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U3-Pad3_ d_xnor		
U4  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U4-Pad3_ d_xnor		
U5  Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U5-Pad3_ d_xnor		
U6  Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U6-Pad3_ d_xnor		
U7  Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U7-Pad3_ d_xnor		
U8  Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U8-Pad3_ d_xnor		
U9  Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U11-Pad1_ d_xnor		
U10  Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U10-Pad3_ d_xnor		
X1  Net-_U3-Pad3_ Net-_U4-Pad3_ Net-_U5-Pad3_ Net-_X1-Pad4_ 3_and		
X2  Net-_U6-Pad3_ Net-_U7-Pad3_ Net-_U8-Pad3_ Net-_X2-Pad4_ 3_and		
U11  Net-_U11-Pad1_ Net-_U10-Pad3_ Net-_U11-Pad3_ d_and		
X3  Net-_U2-Pad2_ Net-_X1-Pad4_ Net-_X2-Pad4_ Net-_U11-Pad3_ Net-_U12-Pad1_ 4_and		
U12  Net-_U12-Pad1_ Net-_U1-Pad18_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U1-Pad18_ PORT		

.end
