* C:\FOSSEE\eSim\library\SubcircuitLibrary\M5234_final\M5234_final.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/12/25 14:19:05

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X2  Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad12_ Net-_U1-Pad1_ Net-_U1-Pad3_ COMPARATOR		
X4  Net-_U1-Pad11_ Net-_U1-Pad10_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad3_ COMPARATOR		
X1  Net-_U1-Pad5_ Net-_U1-Pad4_ Net-_U1-Pad12_ Net-_U1-Pad2_ Net-_U1-Pad3_ COMPARATOR		
X3  Net-_U1-Pad9_ Net-_U1-Pad8_ Net-_U1-Pad12_ Net-_U1-Pad14_ Net-_U1-Pad3_ COMPARATOR		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT		

.end
