* /home/saurabh/Downloads/eSim-1.1.2/Examples/Differentiator/Differentiator.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Mar  8 14:40:54 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R2-Pad2_ Net-_C1-Pad2_ out UA741		
R3  out Net-_C1-Pad2_ 10k		
R1  Net-_C1-Pad1_ in 100k		
R2  GND Net-_R2-Pad2_ 1k		
R4  GND out 1k		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 20n		
v1  in GND pwl		
U1  in plot_v1		
U2  out plot_v1		

.end
