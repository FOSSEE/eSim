* /home/bhargav/eSim-Workspace/IB3858_SPEAKER_CHARACTERISTICS/IB3858_SPEAKER_CHARACTERISTICS.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jul  2 12:52:57 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  v_vr GND SPEAKER		
v1  Net-_R1-Pad1_ GND AC		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 10		
U2  v_vr plot_v1		
U1  Net-_R1-Pad2_ v_vr plot_i2		

.end
