.title KiCad schematic
M2 Net-_M10-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M10-Pad1_ eSim_MOS_P
M1 Net-_M1-Pad1_ Net-_M1-Pad2_ GND GND eSim_MOS_N
U1 Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M3-Pad1_ Net-_M5-Pad2_ Net-_M5-Pad1_ GND Net-_M7-Pad1_ Net-_M7-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad2_ Net-_M11-Pad1_ Net-_M11-Pad2_ Net-_M10-Pad1_ PORT
M8 Net-_M10-Pad1_ Net-_M7-Pad2_ Net-_M7-Pad1_ Net-_M10-Pad1_ eSim_MOS_P
M7 Net-_M7-Pad1_ Net-_M7-Pad2_ GND GND eSim_MOS_N
M5 Net-_M5-Pad1_ Net-_M5-Pad2_ GND GND eSim_MOS_N
M6 Net-_M10-Pad1_ Net-_M5-Pad2_ Net-_M5-Pad1_ Net-_M10-Pad1_ eSim_MOS_P
M10 Net-_M10-Pad1_ Net-_M10-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad1_ eSim_MOS_P
M9 Net-_M10-Pad3_ Net-_M10-Pad2_ GND GND eSim_MOS_N
M12 Net-_M10-Pad1_ Net-_M11-Pad2_ Net-_M11-Pad1_ Net-_M10-Pad1_ eSim_MOS_P
M11 Net-_M11-Pad1_ Net-_M11-Pad2_ GND GND eSim_MOS_N
M3 Net-_M3-Pad1_ Net-_M3-Pad2_ GND GND eSim_MOS_N
M4 Net-_M10-Pad1_ Net-_M3-Pad2_ Net-_M3-Pad1_ Net-_M10-Pad1_ eSim_MOS_P
.end
