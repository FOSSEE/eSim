* C:\FOSSEE\eSim\library\SubcircuitLibrary\Tri_state_buffer\Tri_state_buffer.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/29/25 11:44:13

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M2  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M5  Net-_M5-Pad1_ Net-_M3-Pad2_ Net-_M5-Pad3_ Net-_M1-Pad3_ mosfet_n		
M6  Net-_M5-Pad3_ Net-_M1-Pad1_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_n		
M8  Net-_M5-Pad1_ Net-_M3-Pad1_ Net-_M7-Pad1_ Net-_M2-Pad3_ mosfet_p		
M7  Net-_M7-Pad1_ Net-_M1-Pad1_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_n		
M4  Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M3  Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_n		
U1  Net-_M1-Pad2_ Net-_M3-Pad2_ Net-_M2-Pad3_ Net-_M1-Pad3_ Net-_M5-Pad1_ PORT		

.end
