* C:\FOSSEE\eSim\library\SubcircuitLibrary\AN1186\AN1186.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/10/25 21:13:46

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ d_flop		
U5  Net-_U1-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U3-Pad11_ d_flop		
U7  Net-_U3-Pad11_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U10-Pad1_ d_flop		
U10  Net-_U10-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U10-Pad4_ d_flop		
U2  Net-_U2-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U2-Pad4_ d_flop		
U6  Net-_U6-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U3-Pad6_ d_flop		
U8  Net-_U3-Pad6_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U11-Pad1_ d_flop		
U11  Net-_U11-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U11-Pad4_ d_flop		
U12  Net-_U11-Pad4_ Net-_U12-Pad2_ Net-_U1-Pad1_ d_xor		
U4  Net-_U10-Pad4_ Net-_U1-Pad1_ Net-_U2-Pad1_ d_xor		
U9  Net-_U2-Pad4_ Net-_U1-Pad1_ Net-_U6-Pad1_ d_xor		
U3  Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U12-Pad2_ Net-_U11-Pad4_ Net-_U11-Pad1_ Net-_U3-Pad6_ ? Net-_U2-Pad4_ Net-_U10-Pad4_ Net-_U10-Pad1_ Net-_U3-Pad11_ Net-_U1-Pad4_ ? ? PORT		

.end
