* C:\Users\Shanthipriya\Desktop\madeeasy\FOSSEE\eSim\library\SubcircuitLibrary\74ls90\74ls90.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/15/25 15:54:08

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  /JK /JK /CLK /R01 /R91 /QA ? d_jkff		
U4  Net-_U3-Pad3_ Net-_U3-Pad3_ /CLK /R01 /R91 /QB ? d_jkff		
U8  Net-_U5-Pad3_ Net-_U5-Pad3_ /CLK /R01 /R91 /QC ? d_jkff		
U11  Net-_U10-Pad3_ Net-_U10-Pad3_ /CLK /R01 /R91 /QD Net-_U11-Pad7_ d_jkff		
U3  Net-_U11-Pad7_ /QA Net-_U3-Pad3_ d_and		
U5  /QA /QB Net-_U5-Pad3_ d_and		
U7  /QA /QD Net-_U10-Pad2_ d_and		
U6  /QA /QB Net-_U6-Pad3_ d_and		
U9  Net-_U6-Pad3_ /QC Net-_U10-Pad1_ d_and		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ d_or		
U1  /R91 /CLK /R01 /JK ? ? ? ? /QA /QB /QC /QD PORT		

.end
