.title KiCad schematic
U2 vout plot_v1
X1 unconnected-_X1-Pad1_ vout vin GND unconnected-_X1-Pad5_ vout Net-_X1-Pad7_ unconnected-_X1-Pad8_ LT1007
v3 Net-_X1-Pad7_ GND DC
U1 vin plot_v1
Vv1 vin GND sin(2.5 1.0 1k)
.end
