* E:\IC_CD4037\IC_CD4037.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/17/25 19:14:43

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U6  A Net-_U6-Pad2_ adc_bridge_1		
U7  B Net-_U7-Pad2_ adc_bridge_1		
U8  C1 Net-_U8-Pad2_ adc_bridge_1		
U9  C2 Net-_U9-Pad2_ adc_bridge_1		
U10  C3 Net-_U10-Pad2_ adc_bridge_1		
U11  Net-_U11-Pad1_ D1 dac_bridge_1		
U12  Net-_U12-Pad1_ E1 dac_bridge_1		
U13  Net-_U13-Pad1_ D2 dac_bridge_1		
U14  Net-_U14-Pad1_ E2 dac_bridge_1		
U15  Net-_U15-Pad1_ D3 dac_bridge_1		
U16  Net-_U16-Pad1_ E3 dac_bridge_1		
v1  A GND pulse		
v2  B GND pulse		
v3  C1 GND pulse		
v4  C2 GND pulse		
v5  C3 GND pulse		
U17  D1 plot_v1		
U18  E1 plot_v1		
U19  D2 plot_v1		
U20  E2 plot_v1		
U21  D3 plot_v1		
U22  E3 plot_v1		
U1  A plot_v1		
U2  B plot_v1		
U3  C1 plot_v1		
U4  C2 plot_v1		
U5  C3 plot_v1		
X1  Net-_U8-Pad2_ Net-_U9-Pad2_ Net-_U10-Pad2_ Net-_U7-Pad2_ Net-_U6-Pad2_ Net-_U11-Pad1_ Net-_U12-Pad1_ Net-_U13-Pad1_ Net-_U14-Pad1_ Net-_U15-Pad1_ Net-_U16-Pad1_ CD4037		

.end
