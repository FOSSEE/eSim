* /home/fossee/UpdatedExamples/InvertingAmplifier/InvertingAmplifier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Mar  3 22:37:06 2016

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R4-Pad1_ Net-_R1-Pad2_ out UA741		
R1  in Net-_R1-Pad2_ 1k		
R2  Net-_R1-Pad2_ out 5k		
v1  in GND sine		
R3  out GND 1k		
R4  Net-_R4-Pad1_ GND 1k		
U1  in plot_v1		
U2  out plot_v1		

.end
