* C:\Users\Chaithu\FOSSEE\eSim\library\SubcircuitLibrary\registered_transceiver\registered_transceiver.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 6/7/2025 5:33:15 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U14  Net-_U1-Pad1_ Net-_U1-Pad3_ Net-_U14-Pad3_ d_or		
U12  Net-_U12-Pad1_ Net-_U1-Pad3_ Net-_U12-Pad3_ d_or		
U19  Net-_U19-Pad1_ Net-_U1-Pad5_ Net-_U1-Pad7_ tristate_buff		
U8  Net-_U1-Pad1_ Net-_U12-Pad1_ d_inverter		
U13  Net-_U13-Pad1_ Net-_U13-Pad2_ Net-_U13-Pad3_ d_ff		
U7  Net-_U1-Pad2_ Net-_U12-Pad3_ Net-_U5-Pad1_ d_ff		
U18  Net-_U1-Pad6_ Net-_U1-Pad8_ Net-_U13-Pad2_ d_or		
U20  Net-_U20-Pad1_ Net-_U1-Pad6_ Net-_U20-Pad3_ d_or		
U22  Net-_U1-Pad8_ Net-_U20-Pad1_ d_inverter		
U5  Net-_U5-Pad1_ Net-_U14-Pad3_ Net-_U19-Pad1_ d_ff		
U24  Net-_U1-Pad7_ Net-_U20-Pad3_ Net-_U13-Pad1_ d_ff		
U17  Net-_U13-Pad3_ Net-_U17-Pad2_ Net-_U1-Pad2_ tristate_buff		
U9  Net-_U1-Pad4_ Net-_U17-Pad2_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ PORT		

.end
