* C:\FOSSEE\eSim\library\SubcircuitLibrary\CA3000\CA3000.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 1/4/2026 6:25:27 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
R3  Net-_Q1-Pad1_ Net-_Q2-Pad1_ 8k		
Q2  Net-_Q2-Pad1_ Net-_Q1-Pad3_ Net-_Q2-Pad3_ eSim_NPN		
R1  Net-_Q1-Pad3_ Net-_R1-Pad2_ 4.8k		
R5  Net-_Q2-Pad3_ Net-_Q3-Pad1_ 50		
R9  Net-_Q3-Pad1_ Net-_Q4-Pad3_ 50		
Q4  Net-_Q4-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad3_ eSim_NPN		
R10  Net-_Q1-Pad1_ Net-_Q4-Pad1_ 8k		
Q5  Net-_Q1-Pad1_ Net-_Q5-Pad2_ Net-_Q4-Pad2_ eSim_NPN		
R11  Net-_Q4-Pad2_ Net-_R1-Pad2_ 4.8k		
Q3  Net-_Q3-Pad1_ Net-_Q3-Pad2_ Net-_Q3-Pad3_ eSim_NPN		
R7  Net-_Q3-Pad3_ Net-_R7-Pad2_ 1k		
R4  Net-_Q3-Pad2_ Net-_D1-Pad1_ 2.8k		
R2  Net-_Q3-Pad2_ Net-_R2-Pad2_ 5k		
R8  Net-_R7-Pad2_ Net-_R1-Pad2_ 2k		
R6  Net-_D2-Pad2_ Net-_R1-Pad2_ 2.2k		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
D2  Net-_D1-Pad2_ Net-_D2-Pad2_ eSim_Diode		
U1  Net-_Q1-Pad2_ Net-_R2-Pad2_ Net-_R1-Pad2_ Net-_R7-Pad2_ Net-_D1-Pad1_ Net-_Q5-Pad2_ ? Net-_Q4-Pad1_ Net-_Q1-Pad1_ Net-_Q2-Pad1_ PORT		

.end
