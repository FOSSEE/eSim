* /home/saurabh/Desktop/eSim/Examples/Integrator/Integrator.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Mar 11 16:27:08 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R2-Pad1_ Net-_C1-Pad2_ out UA741		
v1  in GND pwl		
U1  in plot_v1		
U2  out plot_v1		
R1  in Net-_C1-Pad2_ 10k		
R2  Net-_R2-Pad1_ GND 1k		
R3  out Net-_C1-Pad2_ 100k		
C1  out Net-_C1-Pad2_ 100n		
R4  GND out 1k		

.end
