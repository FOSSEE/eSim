* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jun 17 14:53:06 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ D		
D3  Net-_D3-Pad1_ Net-_D1-Pad2_ D		
D4  GND Net-_D3-Pad1_ D		
D2  GND Net-_D1-Pad1_ D		
R1  Net-_D1-Pad2_ GND 1000		
v1  Net-_D1-Pad1_ Net-_D3-Pad1_ sine		

.end
