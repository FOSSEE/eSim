* C:\FOSSEE\eSim\library\SubcircuitLibrary\M5223_My\M5223_My.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/05/25 00:22:44

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q4  Net-_C1-Pad2_ Net-_Q2-Pad1_ Net-_I4-Pad2_ eSim_NPN		
Q2  Net-_Q2-Pad1_ Net-_Q1-Pad3_ Net-_I1-Pad2_ eSim_PNP		
Q1  GND Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_PNP		
Q5  Net-_C1-Pad2_ Net-_Q5-Pad2_ Net-_I1-Pad2_ eSim_PNP		
Q6  GND Net-_Q6-Pad2_ Net-_Q5-Pad2_ eSim_PNP		
Q3  Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_I4-Pad2_ eSim_NPN		
I1  Net-_I1-Pad1_ Net-_I1-Pad2_ dc		
Q11  Net-_I1-Pad1_ Net-_C1-Pad1_ Net-_Q11-Pad3_ eSim_NPN		
Q12  Net-_I1-Pad1_ Net-_Q11-Pad3_ Net-_Q10-Pad2_ eSim_NPN		
Q7  Net-_I4-Pad2_ Net-_C1-Pad2_ Net-_I2-Pad2_ eSim_PNP		
Q8  Net-_I1-Pad1_ Net-_I2-Pad2_ Net-_Q8-Pad3_ eSim_NPN		
Q9  Net-_C1-Pad1_ Net-_Q8-Pad3_ Net-_I4-Pad2_ eSim_NPN		
I2  Net-_I1-Pad1_ Net-_I2-Pad2_ dc		
I3  Net-_I1-Pad1_ Net-_C1-Pad1_ dc		
Q10  Net-_C1-Pad1_ Net-_Q10-Pad2_ Net-_I4-Pad1_ eSim_NPN		
I4  Net-_I4-Pad1_ Net-_I4-Pad2_ dc		
Q13  Net-_I4-Pad2_ Net-_C1-Pad1_ Net-_I4-Pad1_ eSim_PNP		
R3  Net-_Q10-Pad2_ Net-_I4-Pad1_ 500		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 15p		
U1  Net-_Q1-Pad2_ Net-_Q6-Pad2_ Net-_I4-Pad2_ Net-_I1-Pad1_ Net-_I4-Pad1_ PORT		

.end
