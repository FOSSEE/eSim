* C:\FOSSEE\eSim\library\SubcircuitLibrary\tda7050\tda7050.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/08/25 21:45:08

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  ? Net-_U1-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad5_ ? Net-_U1-Pad7_ Net-_U1-Pad8_ ? lm_741		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ PORT		
X2  ? Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad8_ ? Net-_U1-Pad6_ Net-_U1-Pad5_ ? lm_741		

.end
