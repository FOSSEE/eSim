* C:\Users\senba\eSim-Workspace\SN7475_TEST\SN7475_TEST.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/28/25 20:29:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  C D Net-_U3-Pad3_ Net-_U3-Pad4_ adc_bridge_2		
v1  C GND pulse		
v2  D GND pulse		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Q Qbar dac_bridge_2		
U1  C plot_v1		
U2  D plot_v1		
U5  Q plot_v1		
U6  Qbar plot_v1		
X1  Net-_U4-Pad1_ Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U4-Pad2_ SN74LS75		

.end
