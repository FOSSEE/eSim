* C:\FOSSEE\eSim\library\SubcircuitLibrary\74LVC2G00\74LVC2G00.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/16/26 01:20:20

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ CMOS_NAND		
X2  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ CMOS_NAND		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ PORT		

.end
