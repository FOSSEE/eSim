* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/Y9/Y9.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Jul  5 20:37:19 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad7_ Net-_U1-Pad5_ Net-_U1-Pad6_ Y0		
scmode1  SKY130mode		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ PORT		

.end
