* C:\Users\Aditya\eSim-Workspace\LOG_100\LOG_100.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/17/24 18:49:54

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_X1-Pad6_ GND DC		
v2  Net-_X1-Pad9_ GND DC		
U4  OUT plot_db		
U3  OUT plot_v1		
R1  Net-_R1-Pad1_ GND 1000k		
U5  Net-_R3-Pad1_ I2 plot_i2		
U2  Net-_R2-Pad2_ I1 plot_i2		
v3  I1b GND DC		
v4  I2b GND DC		
R3  Net-_R3-Pad1_ I2b 10k		
R2  I1b Net-_R2-Pad2_ 10k		
X1  I1 Net-_R1-Pad1_ ? OUT ? Net-_X1-Pad6_ OUT ? Net-_X1-Pad9_ ? ? ? ? I2 LOG_100		

.end
