.title KiCad schematic
v2 Net-_U3-Pad1_ GND DC
v3 Net-_U3-Pad3_ GND DC
v1 Net-_U1-Pad1_ GND pulse
v4 CLK GND pulse
U5 GND Net-_U5-Pad2_ GND Net-_U5-Pad4_ GND Net-_U5-Pad6_ Net-_U5-Pad7_ Net-_U5-Pad8_ Net-_U5-Pad9_ Net-_U5-Pad10_ Net-_U5-Pad11_ Net-_U5-Pad12_ Net-_U5-Pad13_ Net-_U5-Pad14_ adc_bridge_7
U4 Net-_U4-Pad1_ OUT dac_bridge_1
X1 Net-_U1-Pad2_ Net-_U3-Pad8_ Net-_U3-Pad9_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ Net-_U3-Pad13_ Net-_U3-Pad14_ Net-_U5-Pad8_ Net-_U5-Pad9_ Net-_U5-Pad10_ Net-_U5-Pad11_ Net-_U4-Pad1_ Net-_U5-Pad12_ Net-_U5-Pad13_ Net-_U5-Pad14_ SN54166
v5 Net-_U5-Pad2_ GND DC
v6 Net-_U5-Pad4_ GND DC
v8 Net-_U5-Pad7_ GND DC
v7 Net-_U5-Pad6_ GND pulse
R1 OUT GND 1k
U6 OUT plot_v1
U2 CLK plot_v1
U1 Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_1
U3 Net-_U3-Pad1_ GND Net-_U3-Pad3_ GND GND CLK GND Net-_U3-Pad8_ Net-_U3-Pad9_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ Net-_U3-Pad13_ Net-_U3-Pad14_ adc_bridge_7
.end
