* C:\FOSSEE\eSim\library\SubcircuitLibrary\tff\tff.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/3/2025 3:33:18 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U1-Pad5_ Net-_U2-Pad2_ Net-_U1-Pad7_ Net-_U1-Pad8_ a1 Net-_U3-Pad6_ d_tff		
U1  t clk GND reset Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ adc_bridge_4		
U5  a1 q dac_bridge_1		
U4  Net-_U3-Pad6_ qb dac_bridge_1		
U2  Net-_U1-Pad6_ Net-_U2-Pad2_ d_inverter		

.end
