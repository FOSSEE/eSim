* C:\Users\pavithra\eSim-Workspace\xor_test\xor_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/29/25 12:14:05

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  A GND pulse		
v2  B GND pulse		
U4  J plot_v1		
v9  Net-_X1-Pad14_ GND DC		
U1  A plot_v1		
U2  B plot_v1		
X1  A B J ? ? ? GND ? ? ? ? ? ? Net-_X1-Pad14_ CD4030		

.end
