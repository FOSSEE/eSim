* C:\FOSSEE\eSim\library\SubcircuitLibrary\NAND_GATE_FINAL\NAND_GATE_FINAL.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/12/25 21:44:11

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q2  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
R1  Net-_R1-Pad1_ Net-_Q1-Pad2_ 500		
R2  Net-_R1-Pad1_ Net-_Q3-Pad1_ 60k		
R4  Net-_Q4-Pad1_ Net-_R1-Pad1_ 10k		
Q4  Net-_Q4-Pad1_ Net-_Q3-Pad1_ Net-_D1-Pad1_ eSim_NPN		
Q3  Net-_Q3-Pad1_ Net-_Q1-Pad1_ Net-_Q3-Pad3_ eSim_NPN		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q5  Net-_D1-Pad2_ Net-_Q3-Pad3_ GND eSim_NPN		
R3  Net-_Q3-Pad3_ GND 10k		
U1  Net-_Q1-Pad3_ Net-_Q2-Pad3_ Net-_D1-Pad2_ Net-_R1-Pad1_ PORT		

.end
