* C:\Users\Aditya\eSim-Workspace\Logic_Gates\Logic_Gates.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/28/24 11:42:35

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  A GND pulse		
v2  B GND pulse		
R1  OutA GND 1000k		
X1  A OutA NOT_Gate		
X2  B OutB NOT_Gate		
R2  OutB GND 1000k		
U1  A B OutC XOR_Gate		
R3  OutC GND 1000k		

.end
