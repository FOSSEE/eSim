* C:\FOSSEE\eSim\library\SubcircuitLibrary\74ALS10A\74ALS10A.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/30/26 14:55:34

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X3  Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_X3-Pad3_ CMOS_NAND		
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_X1-Pad3_ CMOS_NAND		
X4  Net-_X3-Pad3_ Net-_U1-Pad7_ Net-_U1-Pad10_ CMOS_NAND		
X5  Net-_X1-Pad3_ Net-_U1-Pad8_ Net-_U1-Pad11_ CMOS_NAND		
X2  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_X2-Pad3_ CMOS_NAND		
X6  Net-_X2-Pad3_ Net-_U1-Pad9_ Net-_U1-Pad12_ CMOS_NAND		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ PORT		

.end
