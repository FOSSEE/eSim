* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/2_in_and/2_in_and.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jul  8 12:32:28 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad3_ Net-_U1-Pad2_ Net-_U1-Pad1_ Net-_X1-Pad4_ Net-_U1-Pad4_ NAND_2		
X2  Net-_X1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad5_ CMOS_INVTR		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ PORT		
scmode1  SKY130mode		

.end
