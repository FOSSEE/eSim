* C:\FOSSEE\eSim\library\SubcircuitLibrary\dm74ls51\dm74ls51.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/03/25 20:46:55

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad1_ Net-_U3-Pad1_ 3_and		
X2  Net-_U1-Pad11_ Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U3-Pad2_ 3_and		
U5  Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U4-Pad1_ d_and		
U2  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U2-Pad3_ d_and		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U1-Pad8_ d_nor		
U4  Net-_U4-Pad1_ Net-_U2-Pad3_ Net-_U1-Pad6_ d_nor		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ PORT		

.end
