* C:\FOSSEE\eSim\library\SubcircuitLibrary\74HC32\74HC32.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/16/2025 7:54:48 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ d_or		
U3  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ d_or		
U4  Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad8_ d_or		
U5  Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad11_ d_or		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ ? Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ ? PORT		

.end
