* /home/saurabh/eSim-Workspace/CMOS_NAND_Gate/CMOS_NAND_Gate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Apr 24 09:28:35 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  inputA GND pulse		
v2  inputB GND pulse		
U2  inputB plot_v1		
U1  inputA plot_v1		
U3  out plot_v1		
X1  inputA inputB out CMOS_NAND		

.end
