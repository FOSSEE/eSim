* E:\IC_SN54H87\IC_SN54H87.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/02/25 10:24:36

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad2_ Net-_U2-Pad2_ Net-_U3-Pad2_ Net-_U4-Pad2_ Net-_U5-Pad2_ Net-_U6-Pad2_ Net-_U9-Pad1_ Net-_U10-Pad1_ Net-_U8-Pad1_ Net-_U7-Pad1_ ? ? ? ? SN54H87		
U1  B Net-_U1-Pad2_ adc_bridge_1		
U2  C Net-_U2-Pad2_ adc_bridge_1		
U3  A1 Net-_U3-Pad2_ adc_bridge_1		
U4  A2 Net-_U4-Pad2_ adc_bridge_1		
U5  A3 Net-_U5-Pad2_ adc_bridge_1		
U6  A4 Net-_U6-Pad2_ adc_bridge_1		
U7  Net-_U7-Pad1_ Y1 dac_bridge_1		
U8  Net-_U8-Pad1_ Y2 dac_bridge_1		
U9  Net-_U9-Pad1_ Y3 dac_bridge_1		
U10  Net-_U10-Pad1_ Y4 dac_bridge_1		
U11  Y1 plot_v1		
U12  Y2 plot_v1		
U13  Y3 plot_v1		
U14  Y4 plot_v1		
v1  B GND pulse		
v2  C GND pulse		
v3  A1 GND pulse		
v4  A2 GND pulse		
v5  A3 GND pulse		
v6  A4 GND pulse		

.end
