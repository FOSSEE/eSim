* C:\Users\Chaithu\FOSSEE\eSim\library\SubcircuitLibrary\SN54HC164\SN54HC164.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/29/2025 7:41:54 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U1-Pad2_ Net-_U1-Pad1_ Net-_U3-Pad1_ d_and		
U2  Net-_U1-Pad3_ Net-_U10-Pad2_ d_buffer		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ PORT		
U7  Net-_U1-Pad5_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad7_ dff_rst		
U3  Net-_U3-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad5_ dff_rst		
U9  Net-_U1-Pad7_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad9_ dff_rst		
U11  Net-_U1-Pad9_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad11_ dff_rst		
U5  Net-_U1-Pad11_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad6_ dff_rst		
U8  Net-_U1-Pad6_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad8_ dff_rst		
U10  Net-_U1-Pad8_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad10_ dff_rst		
U12  Net-_U1-Pad10_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U1-Pad12_ dff_rst		
U6  Net-_U1-Pad4_ Net-_U10-Pad3_ d_inverter		

.end
