.title KiCad schematic
U6 V_Y5 plot_v1
U4 V_Y3 plot_v1
U3 V_Y2 plot_v1
U2 V_Y1 plot_v1
U1 V_Y0 plot_v1
U5 V_Y4 plot_v1
U11 V_Y9 plot_v1
U12 V_Y8 plot_v1
U13 V_Y7 plot_v1
U14 V_D plot_v1
U9 V_A V_B V_C V_D Net-_U9-Pad5_ Net-_U9-Pad6_ Net-_U9-Pad7_ Net-_U9-Pad8_ adc_bridge_4
v1 Net-_X1-Pad16_ GND 5
R7 GND V_Y6 1k
U8 Net-_U8-Pad1_ Net-_U8-Pad2_ Net-_U8-Pad3_ Net-_U8-Pad4_ Net-_U8-Pad5_ Net-_U8-Pad6_ Net-_U8-Pad7_ V_Y0 V_Y1 V_Y2 V_Y3 V_Y4 V_Y5 V_Y6 dac_bridge_7
X1 Net-_U8-Pad1_ Net-_U8-Pad2_ Net-_U8-Pad3_ Net-_U8-Pad4_ Net-_U8-Pad5_ Net-_U8-Pad6_ Net-_U8-Pad7_ GND Net-_U10-Pad3_ Net-_U10-Pad2_ Net-_U10-Pad1_ Net-_U9-Pad8_ Net-_U9-Pad7_ Net-_U9-Pad6_ Net-_U9-Pad5_ Net-_X1-Pad16_ 74145
R5 GND V_Y4 1k
R6 GND V_Y5 1k
R4 GND V_Y3 1k
R1 GND V_Y0 1k
R3 GND V_Y2 1k
R2 GND V_Y1 1k
v_C1 V_C GND DC
R9 GND V_Y8 1k
R8 GND V_Y9 1k
v_B1 V_B GND DC
R10 GND V_Y7 1k
v_D1 V_D GND DC
U10 Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ V_Y9 V_Y8 V_Y7 dac_bridge_3
U17 V_A plot_v1
U16 V_B plot_v1
U15 V_C plot_v1
v_A1 V_A GND DC
U7 V_Y6 plot_v1
.end
