* /home/mallikarjuna/Downloads/eSim-1.1.2/src/SubcircuitLibrary/2bit_upcounter/2bit_upcounter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Jun 22 11:44:38 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U2-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U2-Pad1_ d_dff		
U3  Net-_U3-Pad1_ Net-_U2-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad4_ Net-_U3-Pad1_ d_dff		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ PORT		

.end
