* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jun 24 11:31:48 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U2  1 4 3 d_xor		
U3  1 4 2 d_and		
U1  1 4 3 2 PORT		

.end
