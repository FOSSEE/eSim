* C:\esim\eSim\src\SubcircuitLibrary\Full-Adder\Full-Adder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/21/19 17:15:52

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ PORT		
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad3_ d_xor		
U5  Net-_U2-Pad3_ Net-_U1-Pad3_ Net-_U1-Pad4_ d_xor		
U4  Net-_U2-Pad3_ Net-_U1-Pad3_ Net-_U4-Pad3_ d_and		
U3  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U3-Pad3_ d_and		
U6  Net-_U3-Pad3_ Net-_U4-Pad3_ Net-_U1-Pad5_ d_or		

.end
