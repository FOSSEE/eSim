* E:\FOSSEE\eSim\library\SubcircuitLibrary\HEF4531B\HEF4531B.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/24/25 11:35:39

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad3_ d_xor		
U3  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U3-Pad3_ d_xor		
U4  Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U10-Pad1_ d_xor		
U5  Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U10-Pad2_ d_xor		
U6  Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U6-Pad3_ d_xor		
U7  Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U7-Pad3_ d_xor		
U9  Net-_U2-Pad3_ Net-_U3-Pad3_ Net-_U11-Pad1_ d_xor		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ d_xor		
U8  Net-_U6-Pad3_ Net-_U7-Pad3_ Net-_U12-Pad1_ d_xor		
U11  Net-_U11-Pad1_ Net-_U10-Pad3_ Net-_U11-Pad3_ d_xor		
U12  Net-_U12-Pad1_ Net-_U1-Pad13_ Net-_U12-Pad3_ d_xor		
U13  Net-_U11-Pad3_ Net-_U12-Pad3_ Net-_U13-Pad3_ d_xor		
U14  Net-_U13-Pad3_ Net-_U1-Pad16_ d_buffer		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ ? ? Net-_U1-Pad16_ PORT		

.end
