* /home/bhargav/Downloads/eSim-1.1.2/src/SubcircuitLibrary/LM3046/LM3046.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Jun 22 11:57:18 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
Q4  Net-_Q4-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad3_ eSim_NPN		
Q5  Net-_Q5-Pad1_ Net-_Q5-Pad2_ Net-_Q5-Pad3_ eSim_NPN		
Q3  Net-_Q3-Pad1_ Net-_Q3-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
U1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ Net-_Q3-Pad2_ Net-_Q3-Pad1_ Net-_Q5-Pad2_ Net-_Q5-Pad3_ Net-_Q5-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad3_ Net-_Q4-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ Net-_Q2-Pad1_ PORT		

.end
