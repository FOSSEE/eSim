* D:\FOSSEE\eSim\library\SubcircuitLibrary\SN74177\SN74177.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/13/25 09:20:10

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U6  Net-_U16-Pad3_ Net-_U14-Pad2_ Net-_U6-Pad3_ d_nand		
U7  Net-_U17-Pad3_ Net-_U14-Pad2_ Net-_U7-Pad3_ d_nand		
U8  Net-_U19-Pad3_ Net-_U14-Pad2_ Net-_U8-Pad3_ d_nand		
U9  Net-_U18-Pad3_ Net-_U14-Pad2_ Net-_U9-Pad3_ d_nand		
U2  /13 Net-_U16-Pad2_ d_buffer		
U3  /1 /13 Net-_U14-Pad2_ d_nand		
U1  /1 /2 /3 /4 /5 /6 ? /8 /9 /10 /11 /12 /13 ? PORT		
U4  /4 Net-_U14-Pad2_ Net-_U16-Pad1_ d_and		
U16  Net-_U16-Pad1_ Net-_U16-Pad2_ Net-_U16-Pad3_ d_nand		
U5  /10 Net-_U14-Pad2_ Net-_U17-Pad1_ d_and		
U17  Net-_U17-Pad1_ Net-_U16-Pad2_ Net-_U17-Pad3_ d_nand		
U15  /3 Net-_U14-Pad2_ Net-_U15-Pad3_ d_and		
U19  Net-_U15-Pad3_ Net-_U16-Pad2_ Net-_U19-Pad3_ d_nand		
U14  /11 Net-_U14-Pad2_ Net-_U14-Pad3_ d_and		
U18  Net-_U14-Pad3_ Net-_U16-Pad2_ Net-_U18-Pad3_ d_nand		
X1  ? /8 Net-_U6-Pad3_ ? /5 Net-_U16-Pad3_ tff_1		
X4  ? /2 Net-_U9-Pad3_ ? /12 Net-_U18-Pad3_ tff_1		
X3  ? /9 Net-_U8-Pad3_ ? /2 Net-_U19-Pad3_ tff_1		
X2  ? /6 Net-_U7-Pad3_ ? /9 Net-_U17-Pad3_ tff_1		

.end
