* C:\FOSSEE\eSim\library\SubcircuitLibrary\74LS90\74LS90.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/24/25 17:57:37

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U7  ? ? Net-_U5-Pad2_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U7-Pad6_ ? d_jkff		
U12  ? ? Net-_U10-Pad6_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U12-Pad6_ ? d_jkff		
U10  Net-_U10-Pad1_ ? Net-_U10-Pad3_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U10-Pad6_ ? d_jkff		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U10-Pad5_ d_nand		
U6  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U10-Pad4_ d_nand		
U15  Net-_U14-Pad3_ Net-_U15-Pad2_ Net-_U10-Pad3_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U15-Pad2_ Net-_U10-Pad1_ d_srff		
U5  Net-_U1-Pad1_ Net-_U5-Pad2_ adc_bridge_1		
U8  Net-_U1-Pad6_ Net-_U10-Pad3_ adc_bridge_1		
U14  Net-_U10-Pad6_ Net-_U12-Pad6_ Net-_U14-Pad3_ d_and		
U2  Net-_U1-Pad2_ Net-_U1-Pad4_ Net-_U2-Pad3_ Net-_U2-Pad4_ adc_bridge_2		
U4  Net-_U1-Pad3_ Net-_U1-Pad5_ Net-_U3-Pad1_ Net-_U3-Pad2_ adc_bridge_2		
U9  Net-_U7-Pad6_ Net-_U1-Pad7_ dac_bridge_1		
U11  Net-_U10-Pad6_ Net-_U1-Pad8_ dac_bridge_1		
U16  Net-_U15-Pad2_ Net-_U1-Pad10_ dac_bridge_1		
U13  Net-_U12-Pad6_ Net-_U1-Pad9_ dac_bridge_1		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ PORT		

.end
