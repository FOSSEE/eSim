* eeschema netlist version 1.1 (spice format) creation date: monday 17 december 2012 10:57:49 am ist

* Inverter d_inverter
* SR Latch d_srlatch
e2  18 0 23 14 10000
* Limiter limit8
* Digital to Analog converter dac8
* Analog to Digital converter adc8
u1  22 14 7 6 15 16 3 13 port
r8  9 2 1500
q1 3 2 22 qnom
r7  18 20 25
r6  17 19 25
e1  17 0 16 15 10000
r4  16 15 2e6
r5  23 14 2e6
r3  23 22 5000
r2  15 23 5000
r1  13 15 5000
a1 5 21 u5
.model u5 d_inverter(rise_delay=1e-12 fall_delay=1e-12 input_load=1e-12)
a2 1 4 5 21 21 8 10 u6
.model u6 d_srlatch(rise_delay=1e-12 fall_delay=1e-12 ic=0
+sr_load=1e-12 enable_load=1e-12 set_load=1e-12 reset_load=1e-12
+sr_delay=1e-12 enable_delay=1e-12 set_delay=1e-12 reset_delay=1e-12)
a3 19 11 u4
a4 20 12 u4
.model u4 limit(out_lower_limit=0.0 out_upper_limit=5.0)
a5 [8] [7] u3
a6 [10] [9] u3
.model u3 dac_bridge(out_low=0.2 out_high=5.0 out_undef=5.0 )
a7 [11] [4] u2
a8 [12] [1] u2
a9 [6] [5] u2
.model u2 adc_bridge(in_low=0.8 in_high=2.0 )
