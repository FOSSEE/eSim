.title KiCad schematic
U8 Net-_U10-Pad1_ Net-_U8-Pad2_ Net-_U15-Pad1_ d_and
U7 Net-_U11-Pad1_ Net-_U7-Pad2_ Net-_U14-Pad2_ d_and
U6 Net-_U10-Pad1_ Net-_U6-Pad2_ Net-_U14-Pad1_ d_and
U10 Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ d_and
U9 Net-_U11-Pad1_ Net-_U9-Pad2_ Net-_U15-Pad2_ d_and
U5 Net-_U4-Pad1_ Net-_U11-Pad1_ d_buffer
U3 Net-_U3-Pad1_ Net-_U18-Pad2_ d_inverter
U4 Net-_U4-Pad1_ Net-_U10-Pad1_ d_inverter
U1 Net-_U4-Pad1_ Net-_U6-Pad2_ Net-_U7-Pad2_ Net-_U18-Pad3_ Net-_U8-Pad2_ Net-_U9-Pad2_ Net-_U19-Pad3_ unconnected-_U1-Pad8_ Net-_U20-Pad3_ Net-_U11-Pad2_ Net-_U10-Pad2_ Net-_U21-Pad3_ Net-_U13-Pad2_ Net-_U12-Pad2_ Net-_U3-Pad1_ unconnected-_U1-Pad16_ PORT
U17 Net-_U12-Pad3_ Net-_U13-Pad3_ Net-_U17-Pad3_ d_or
U16 Net-_U10-Pad3_ Net-_U11-Pad3_ Net-_U16-Pad3_ d_or
U15 Net-_U15-Pad1_ Net-_U15-Pad2_ Net-_U15-Pad3_ d_or
U19 Net-_U15-Pad3_ Net-_U18-Pad2_ Net-_U19-Pad3_ d_tristate
U21 Net-_U17-Pad3_ Net-_U18-Pad2_ Net-_U21-Pad3_ d_tristate
U20 Net-_U16-Pad3_ Net-_U18-Pad2_ Net-_U20-Pad3_ d_tristate
U18 Net-_U14-Pad3_ Net-_U18-Pad2_ Net-_U18-Pad3_ d_tristate
U14 Net-_U14-Pad1_ Net-_U14-Pad2_ Net-_U14-Pad3_ d_or
U13 Net-_U11-Pad1_ Net-_U13-Pad2_ Net-_U13-Pad3_ d_and
U12 Net-_U10-Pad1_ Net-_U12-Pad2_ Net-_U12-Pad3_ d_and
U11 Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ d_and
.end
