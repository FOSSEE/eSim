* C:\FOSSEE\eSim\library\SubcircuitLibrary\74HC125\74HC125.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/16/2025 10:09:01 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U1-Pad3_ Net-_U2-Pad2_ Net-_U1-Pad5_ d_tristate		
U5  Net-_U1-Pad4_ Net-_U3-Pad2_ Net-_U1-Pad6_ d_tristate		
U8  Net-_U1-Pad11_ Net-_U6-Pad2_ Net-_U1-Pad8_ d_tristate		
U9  Net-_U1-Pad12_ Net-_U7-Pad2_ Net-_U1-Pad10_ d_tristate		
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ PORT		
U3  Net-_U1-Pad2_ Net-_U3-Pad2_ d_inverter		
U6  Net-_U1-Pad7_ Net-_U6-Pad2_ d_inverter		
U7  Net-_U1-Pad9_ Net-_U7-Pad2_ d_inverter		

.end
