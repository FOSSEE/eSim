* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/Quad_D_FF/Quad_D_FF.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jun 24 11:58:14 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad8_ D_FF		
X2  Net-_U1-Pad3_ Net-_U1-Pad2_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad9_ D_FF		
X3  Net-_U1-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad10_ D_FF		
X4  Net-_U1-Pad5_ Net-_U1-Pad2_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad11_ D_FF		
X5  Net-_U1-Pad8_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad12_ CMOS_INVTR		
X6  Net-_U1-Pad9_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad13_ CMOS_INVTR		
X7  Net-_U1-Pad10_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad14_ CMOS_INVTR		
X8  Net-_U1-Pad11_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad15_ CMOS_INVTR		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ PORT		
scmode1  SKY130mode		

.end
