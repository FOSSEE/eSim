* C:\FOSSEE\eSim\library\SubcircuitLibrary\CD4010BQ1\CD4010BQ1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/19/25 10:33:51

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad7_ VCC VDD GND 1_CD4010B		
X2  Net-_U1-Pad2_ Net-_U1-Pad8_ VCC VDD GND 1_CD4010B		
X3  Net-_U1-Pad3_ Net-_U1-Pad9_ VCC VDD GND 1_CD4010B		
X4  Net-_U1-Pad4_ Net-_U1-Pad10_ VCC VDD GND 1_CD4010B		
X5  Net-_U1-Pad5_ Net-_U1-Pad11_ VCC VDD GND 1_CD4010B		
X6  Net-_U1-Pad6_ Net-_U1-Pad12_ VCC VDD GND 1_CD4010B		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ VCC VDD GND PORT		

.end
