* eeschema netlist version 1.1 (spice format) creation date: 08/21/14 11:07:22
.include diode.lib

u2  5 8 1 port
* f2
* Analog Switch analogswitch
d1  4 2 diode
v2  3 4 dc 0
c1  5 6 10u
r2  5 6 1
* f1
v1  9 7 dc 0
r1  8 9 50
Vf2 2 5 0
f2 5 6 Vf2 100
Vf1 7 5 0
f1 5 6 Vf1 10
a1 6 (1 3) u1
.model u1 aswitch(cntl_on=0.25 cntl_off=0.1 r_on=0.0125 r_off=1000000)
