* C:\FOSSEE\eSim\library\SubcircuitLibrary\LH0004\LH0004.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/05/25 11:43:58

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_PNP		
Q3  Net-_Q2-Pad3_ Net-_Q1-Pad1_ Net-_Q1-Pad2_ eSim_PNP		
R3  Net-_Q1-Pad3_ Net-_Q1-Pad2_ 40K		
R1  Net-_Q1-Pad1_ Net-_R1-Pad2_ 600K		
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_PNP		
Q4  Net-_Q4-Pad1_ Net-_Q4-Pad2_ Net-_Q2-Pad3_ eSim_PNP		
R2  Net-_Q2-Pad1_ Net-_Q10-Pad1_ 300K		
R4  Net-_Q4-Pad1_ Net-_Q10-Pad1_ 300K		
R5  Net-_Q1-Pad3_ Net-_Q6-Pad3_ 50K		
Q6  Net-_Q5-Pad1_ Net-_Q5-Pad1_ Net-_Q6-Pad3_ eSim_PNP		
Q7  Net-_Q10-Pad2_ Net-_Q5-Pad1_ Net-_Q7-Pad3_ eSim_PNP		
R7  Net-_Q1-Pad3_ Net-_Q7-Pad3_ 50K		
Q5  Net-_Q5-Pad1_ Net-_Q4-Pad1_ Net-_Q5-Pad3_ eSim_NPN		
Q8  Net-_Q10-Pad2_ Net-_Q2-Pad1_ Net-_Q5-Pad3_ eSim_NPN		
R6  Net-_Q5-Pad3_ Net-_Q10-Pad1_ 50K		
Q9  Net-_Q1-Pad3_ Net-_Q10-Pad2_ Net-_Q10-Pad3_ eSim_NPN		
Q10  Net-_Q10-Pad1_ Net-_Q10-Pad2_ Net-_Q10-Pad3_ eSim_PNP		
U1  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q10-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad1_ Net-_Q1-Pad1_ Net-_R1-Pad2_ Net-_Q10-Pad3_ Net-_Q1-Pad3_ Net-_Q10-Pad2_ PORT		

.end
