* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/SN54L99/SN54L99.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Jul 10 18:58:06 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
scmode1  SKY130mode		
X4  Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_X4-Pad3_ Net-_U1-Pad4_ /mode Net-_X1-Pad4_ Net-_U1-Pad13_ Net-_U1-Pad15_ Net-_U1-Pad5_ SerialParallel_blk		
X6  Net-_U1-Pad5_ Net-_X1-Pad4_ /mode Net-_U1-Pad8_ Net-_X4-Pad3_ Net-_U1-Pad13_ Net-_U1-Pad15_ Net-_U1-Pad9_ DS_blk		
X7  Net-_U1-Pad9_ Net-_X1-Pad4_ /mode Net-_U1-Pad10_ Net-_X4-Pad3_ Net-_U1-Pad13_ Net-_U1-Pad15_ Net-_U1-Pad11_ DS_blk		
X8  Net-_U1-Pad11_ Net-_X1-Pad4_ /mode Net-_U1-Pad12_ Net-_X4-Pad3_ Net-_U1-Pad13_ Net-_U1-Pad15_ Net-_U1-Pad14_ DS_blk		
X2  Net-_U1-Pad13_ Net-_X1-Pad4_ /RS Net-_U1-Pad15_ Net-_X2-Pad5_ 2_in_and		
X3  Net-_U1-Pad13_ /mode /LS Net-_U1-Pad15_ Net-_X3-Pad5_ 2_in_and		
X5  Net-_X2-Pad5_ Net-_X3-Pad5_ Net-_U1-Pad13_ Net-_U1-Pad15_ Net-_X4-Pad3_ or_2		
X1  /mode Net-_U1-Pad13_ Net-_U1-Pad15_ Net-_X1-Pad4_ CMOS_INVTR		
U1  /RS /mode /LS Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ PORT		

.end
