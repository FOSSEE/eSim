* analysis type *
.tran 1n 100n
*
* input sources *
v1 100 0 DC PWL ( 0n 0.0 5n 0.0 5.1n 2.0 10n 0.0 10.1n 2.0 15n 2.0 15.1n 2.0 20n 0 20.1n 2.0 25n 2.0 25.1n 2.0 30n 2.0 30.1n 2.0
               + 40n 0.0 50n 0.0 50.1n 2.0 60n 2.0 60.1n 0.0 70n 0.0 70.1n 2.0 80n 2.0 80.1n 0.0 90n 0.0 100n 2.0)

v2 200 0 DC PWL ( 0n 2.0 5n 2.0 5.1n 0.0 10n 0.0 10.1n 2.0 15n 2.0 15.1n 0.0 20n 0 20.1n 2.0 25n 2.0 25.1n 0.0 30n 2.0 30.1n 2.0
               + 40n 0.0 50n 0.0 50.1n 2.0 60n 2.0 60.1n 0.0 70n 0.0 70.1n 2.0 80n 2.0 80.1n 0.0 90n 0.0 100n 2.0)

* resistors to ground *
r1 100 0 1k
r2 200 0 1k

rload1 300 0 10k
rload2 400 0 10k
*
* adc_bridge blocks *
aconverter1 [100 200]  [1 2] adc_bridge1

.model adc_bridge1 adc_bridge ( in_low =0.3 in_high =0.7
+ rise_delay =1.0e-12 fall_delay =1.0e-12)

ainverter [1 2] [10 20]  inv1

.model inv1 inverter(instance_id = 101 rise_delay = 1.0e-12 fall_delay = 1.0e-12 stop_time=90e-9)


aconverter2 [10 20] [30 40] dac_bridge1

.model dac_bridge1 dac_bridge( out_low=0.25 out_high=5.0 
+out_undef=1.8 t_rise=0.5e-9 t_fall=0.5e-9) 

.end
 

