* C:\FOSSEE\eSim\library\SubcircuitLibrary\SN74LS00\SN74LS00.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/12/25 21:31:58

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad14_ Nand_gate_final		
X3  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad14_ Nand_gate_final		
X2  Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U1-Pad8_ Net-_U1-Pad14_ Nand_gate_final		
X4  Net-_U1-Pad13_ Net-_U1-Pad12_ Net-_U1-Pad11_ Net-_U1-Pad14_ Nand_gate_final		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ ? Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT		

.end
