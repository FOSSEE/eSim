.title KiCad schematic
U1 Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ unconnected-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ unconnected-_U1-Pad16_ PORT
U20 Net-_U14-Pad3_ Net-_U17-Pad2_ Net-_U1-Pad12_ d_tristate
U13 Net-_U13-Pad1_ Net-_U13-Pad2_ Net-_U13-Pad3_ d_or
U15 Net-_U11-Pad3_ Net-_U12-Pad3_ Net-_U15-Pad3_ d_or
U16 Net-_U16-Pad1_ Net-_U16-Pad2_ Net-_U16-Pad3_ d_or
U19 Net-_U16-Pad3_ Net-_U17-Pad2_ Net-_U1-Pad9_ d_tristate
U14 Net-_U14-Pad1_ Net-_U10-Pad3_ Net-_U14-Pad3_ d_or
U17 Net-_U13-Pad3_ Net-_U17-Pad2_ Net-_U1-Pad7_ d_tristate
U18 Net-_U15-Pad3_ Net-_U17-Pad2_ Net-_U1-Pad4_ d_tristate
U8 Net-_U10-Pad1_ Net-_U1-Pad11_ Net-_U16-Pad2_ d_and
U7 Net-_U11-Pad1_ Net-_U1-Pad10_ Net-_U16-Pad1_ d_and
U11 Net-_U11-Pad1_ Net-_U1-Pad3_ Net-_U11-Pad3_ d_and
U12 Net-_U10-Pad1_ Net-_U1-Pad2_ Net-_U12-Pad3_ d_and
U9 Net-_U11-Pad1_ Net-_U1-Pad13_ Net-_U14-Pad1_ d_and
U10 Net-_U10-Pad1_ Net-_U1-Pad14_ Net-_U10-Pad3_ d_and
U6 Net-_U10-Pad1_ Net-_U1-Pad5_ Net-_U13-Pad2_ d_and
U5 Net-_U11-Pad1_ Net-_U1-Pad6_ Net-_U13-Pad1_ d_and
U3 Net-_U1-Pad15_ Net-_U17-Pad2_ d_inverter
U4 Net-_U10-Pad1_ Net-_U11-Pad1_ d_inverter
U2 Net-_U1-Pad1_ Net-_U10-Pad1_ d_inverter
.end
