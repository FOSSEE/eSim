* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/CD4044BMS/CD4044BMS.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Jun 14 11:29:04 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad11_ Net-_U1-Pad2_ Net-_U1-Pad10_ Net-_U1-Pad1_ Net-_U1-Pad3_ Net-_U1-Pad12_ SR_Latch_with_Enable		
X3  Net-_U1-Pad11_ Net-_U1-Pad2_ Net-_U1-Pad10_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad14_ SR_Latch_with_Enable		
X2  Net-_U1-Pad11_ Net-_U1-Pad2_ Net-_U1-Pad10_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad13_ SR_Latch_with_Enable		
X4  Net-_U1-Pad11_ Net-_U1-Pad2_ Net-_U1-Pad10_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad15_ SR_Latch_with_Enable		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ PORT		
scmode1  SKY130mode		

.end
