* C:\FOSSEE\eSim\library\SubcircuitLibrary\SN54LVC157A\SN54LVC157A.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/23/25 15:20:18

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U9  Net-_U1-Pad4_ Net-_U11-Pad2_ Net-_U16-Pad1_ d_and		
U10  Net-_U1-Pad5_ Net-_U10-Pad2_ Net-_U10-Pad3_ d_and		
U16  Net-_U16-Pad1_ Net-_U10-Pad3_ Net-_U1-Pad6_ d_or		
U11  Net-_U1-Pad7_ Net-_U11-Pad2_ Net-_U11-Pad3_ d_and		
U12  Net-_U1-Pad8_ Net-_U10-Pad2_ Net-_U12-Pad3_ d_and		
U17  Net-_U11-Pad3_ Net-_U12-Pad3_ Net-_U1-Pad9_ d_or		
U13  Net-_U1-Pad10_ Net-_U11-Pad2_ Net-_U13-Pad3_ d_and		
U14  Net-_U1-Pad11_ Net-_U10-Pad2_ Net-_U14-Pad3_ d_and		
U18  Net-_U13-Pad3_ Net-_U14-Pad3_ Net-_U1-Pad12_ d_or		
U7  Net-_U1-Pad1_ Net-_U11-Pad2_ Net-_U15-Pad1_ d_and		
U8  Net-_U1-Pad2_ Net-_U10-Pad2_ Net-_U15-Pad2_ d_and		
U15  Net-_U15-Pad1_ Net-_U15-Pad2_ Net-_U1-Pad3_ d_or		
U5  Net-_U2-Pad2_ Net-_U3-Pad2_ Net-_U11-Pad2_ d_and		
U6  Net-_U4-Pad2_ Net-_U1-Pad14_ Net-_U10-Pad2_ d_and		
U2  Net-_U1-Pad13_ Net-_U2-Pad2_ d_inverter		
U3  Net-_U1-Pad14_ Net-_U3-Pad2_ d_inverter		
U4  Net-_U1-Pad13_ Net-_U4-Pad2_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT		

.end
