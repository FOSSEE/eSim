* C:\FOSSEE\eSim\library\SubcircuitLibrary\CD4040\CD4040.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/3/2025 3:49:12 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  vdd clk q1 rst tff		
X2  vdd q1 q2 rst tff		
X3  vdd q2 q3 rst tff		
X4  vdd q3 q4 rst tff		
X5  vdd q4 q5 rst tff		
X6  vdd q5 q6 rst tff		
X7  vdd q6 q7 rst tff		
X8  vdd q7 q8 rst tff		
X9  vdd q8 q9 rst tff		
X10  vdd q9 q10 rst tff		
X11  vdd q10 q11 rst tff		
X12  vdd q11 q12 rst tff		
v1  vdd GND 5v		

.end
