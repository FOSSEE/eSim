* C:\Users\HP\OneDrive\Documents\FOSSEE\eSim\library\SubcircuitLibrary\ICL7660\ICL7660.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/26/25 17:20:02

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
C1  /Vin /CAP+ 100u		
D1  /CAP+ GND eSim_Diode		
D2  /OUT /CAP+ eSim_Diode		
C2  /OUT GND 100u		
U1  ? /CAP+ GND GND GND /Vin ? /OUT PORT		

.end
