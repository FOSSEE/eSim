* C:\Users\Chaithu\FOSSEE\eSim\library\SubcircuitLibrary\registered_transciever\registered_transciever.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 6/9/2025 2:16:21 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U5-Pad3_ d_or		
U4  Net-_U3-Pad2_ Net-_U1-Pad4_ Net-_U2-Pad2_ d_or		
U3  Net-_U1-Pad3_ Net-_U3-Pad2_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ PORT		
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ d_ff		
U6  Net-_U2-Pad3_ Net-_U5-Pad3_ Net-_U6-Pad3_ d_ff		
U7  Net-_U6-Pad3_ Net-_U1-Pad2_ Net-_U1-Pad5_ tristate_buff		
U10  Net-_U1-Pad8_ Net-_U1-Pad7_ Net-_U10-Pad3_ d_or		
U11  Net-_U11-Pad1_ Net-_U1-Pad7_ Net-_U11-Pad3_ d_or		
U12  Net-_U1-Pad8_ Net-_U11-Pad1_ d_inverter		
U13  Net-_U1-Pad5_ Net-_U11-Pad3_ Net-_U13-Pad3_ d_ff		
U9  Net-_U13-Pad3_ Net-_U10-Pad3_ Net-_U8-Pad1_ d_ff		
U8  Net-_U8-Pad1_ Net-_U1-Pad6_ Net-_U1-Pad1_ tristate_buff		

.end
