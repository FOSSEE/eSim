* C:\FOSSEE\eSim\library\SubcircuitLibrary\74HC157\74HC157.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/10/2025 5:51:02 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad9_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U3-Pad1_ mux		
X2  Net-_U1-Pad9_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U4-Pad1_ mux		
X3  Net-_U1-Pad9_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U5-Pad1_ mux		
X4  Net-_U1-Pad9_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U6-Pad1_ mux		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT		
U3  Net-_U3-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad11_ d_and		
U4  Net-_U4-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad12_ d_and		
U5  Net-_U5-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad13_ d_and		
U6  Net-_U6-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad14_ d_and		
U2  Net-_U1-Pad10_ Net-_U2-Pad2_ d_inverter		

.end
