* C:\FOSSEE\eSim\library\SubcircuitLibrary\3_nor\3_nor.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/13/25 12:25:06

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_n		
M5  Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_n		
M6  Net-_M1-Pad1_ Net-_M4-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_n		
M2  Net-_M2-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad1_ eSim_MOS_P		
M3  Net-_M2-Pad3_ Net-_M3-Pad2_ Net-_M3-Pad3_ Net-_M2-Pad1_ eSim_MOS_P		
M4  Net-_M3-Pad3_ Net-_M4-Pad2_ Net-_M1-Pad1_ Net-_M2-Pad1_ eSim_MOS_P		
U4  Net-_U3-Pad2_ Net-_U1-Pad6_ d_buffer		
U3  Net-_M1-Pad1_ Net-_U3-Pad2_ adc_bridge_1		
U2  Net-_U1-Pad3_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_M1-Pad2_ Net-_M3-Pad2_ Net-_M4-Pad2_ dac_bridge_3		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_M2-Pad1_ Net-_M1-Pad3_ Net-_U1-Pad6_ PORT		

.end
