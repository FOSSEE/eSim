* /home/saurabh/eSim-Workspace/Cmosinvertor/Cmosinvertor.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Nov 27 14:17:36 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  out1 plot_v1		
X1  out7 out1 INVCMOS		
X2  out1 out2 INVCMOS		
X3  out2 out3 INVCMOS		
U3  out2 plot_v1		
U4  out3 plot_v1		
X4  out3 out4 INVCMOS		
U5  out4 plot_v1		
X5  out4 out5 INVCMOS		
U6  out5 plot_v1		
X6  out5 out6 INVCMOS		
U7  out6 plot_v1		
U8  out7 plot_v1		
U9  out6 Net-_U1-Pad1_ adc_bridge_1		
U10  Net-_U1-Pad2_ out7 dac_bridge_1		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ inverter		

.end
