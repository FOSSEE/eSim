* E:\FOSSEE\eSim\library\SubcircuitLibrary\TL560C\TL560C.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/13/25 11:09:02

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
Q3  Net-_Q3-Pad1_ Net-_Q3-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
R1  Net-_Q1-Pad3_ Net-_Q6-Pad3_ 5k		
Q2  Net-_Q2-Pad1_ Net-_Q1-Pad1_ Net-_Q2-Pad3_ eSim_PNP		
Q4  Net-_Q4-Pad1_ Net-_Q3-Pad1_ Net-_Q2-Pad3_ eSim_PNP		
R2  Net-_Q6-Pad2_ Net-_Q2-Pad1_ 1.3k		
Q6  Net-_Q3-Pad2_ Net-_Q6-Pad2_ Net-_Q6-Pad3_ eSim_NPN		
Q5  Net-_Q5-Pad1_ Net-_Q4-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
R3  Net-_R3-Pad1_ Net-_Q3-Pad2_ 2.5k		
R5  Net-_Q6-Pad3_ Net-_R3-Pad1_ 3k		
R4  Net-_R3-Pad1_ Net-_Q2-Pad3_ 1.7k		
Q7  Net-_Q7-Pad1_ Net-_Q5-Pad1_ Net-_Q2-Pad3_ eSim_PNP		
R6  Net-_Q8-Pad1_ Net-_Q2-Pad3_ 0.3k		
Q8  Net-_Q8-Pad1_ Net-_Q7-Pad1_ Net-_Q8-Pad3_ eSim_NPN		
R7  Net-_Q9-Pad2_ Net-_Q8-Pad3_ 0.2k		
Q9  Net-_Q9-Pad1_ Net-_Q9-Pad2_ Net-_Q6-Pad3_ eSim_NPN		
R8  Net-_Q6-Pad3_ Net-_Q9-Pad2_ 3k		
U1  Net-_Q1-Pad2_ Net-_Q2-Pad3_ Net-_Q6-Pad3_ Net-_R3-Pad1_ Net-_Q9-Pad1_ PORT		

.end
