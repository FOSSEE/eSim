* C:\FOSSEE\eSim\library\SubcircuitLibrary\CD4066B\CD4066B.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/09/25 14:21:31

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U2-Pad2_ Net-_U3-Pad2_ d_inverter		
U4  Net-_U3-Pad2_ Net-_U4-Pad2_ d_inverter		
U7  Net-_U4-Pad2_ Net-_U6-Pad1_ d_inverter		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ ? eSim_MOS_P		
M3  Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ ? eSim_MOS_N		
M2  Net-_M1-Pad3_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ eSim_MOS_N		
M4  Net-_M4-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ ? eSim_MOS_P		
M5  Net-_M4-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad1_ Net-_M1-Pad3_ eSim_MOS_N		
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ adc_bridge_1		
U6  Net-_U6-Pad1_ Net-_M1-Pad2_ dac_bridge_1		
U5  Net-_U4-Pad2_ Net-_M3-Pad2_ dac_bridge_1		
U1  Net-_U1-Pad1_ Net-_M1-Pad1_ Net-_M2-Pad3_ Net-_M4-Pad1_ GND PORT		

.end
