* C:\FOSSEE\eSim\library\SubcircuitLibrary\LM431\LM431.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 12/15/24 01:48:32

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  Net-_Q1-Pad3_ Net-_Q2-Pad1_ 12k		
R2  Net-_Q2-Pad2_ Net-_Q2-Pad1_ 800		
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
R3  Net-_Q1-Pad3_ Net-_Q3-Pad1_ 12k		
Q3  Net-_Q3-Pad1_ Net-_Q2-Pad1_ Net-_Q3-Pad3_ eSim_NPN		
R4  Net-_Q3-Pad3_ Net-_Q2-Pad3_ 640		
R5  Net-_Q3-Pad1_ Net-_C1-Pad1_ 2.5k		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 0.1nF		
Q4  Net-_C1-Pad2_ Net-_C1-Pad1_ Net-_Q2-Pad3_ eSim_NPN		
Q5  Net-_C1-Pad2_ Net-_C1-Pad2_ Net-_C2-Pad1_ eSim_PNP		
C2  Net-_C2-Pad1_ Net-_C2-Pad2_ 0.1nF		
Q6  Net-_C2-Pad1_ Net-_C2-Pad2_ Net-_Q6-Pad3_ eSim_NPN		
R6  Net-_Q6-Pad3_ Net-_Q2-Pad3_ 1k		
Q7  Net-_C2-Pad1_ Net-_Q6-Pad3_ Net-_Q7-Pad3_ eSim_NPN		
R7  Net-_Q7-Pad3_ Net-_Q2-Pad3_ 3.3		
Q1  Net-_C2-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
U1  Net-_Q1-Pad2_ Net-_C2-Pad1_ Net-_Q2-Pad3_ PORT		
Q8  Net-_C2-Pad2_ Net-_C1-Pad2_ Net-_C2-Pad1_ eSim_PNP		

.end
