* C:\Users\Aditya\eSim-Workspace\MPY100\MPY100.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/27/24 22:47:08

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_X1-Pad10_ GND DC		
v4  Net-_X1-Pad3_ GND DC		
R2  Net-_R1-Pad2_ Vout 70k		
R1  GND Net-_R1-Pad2_ 10k		
v2  V1 GND sine		
v3  V2 GND sine		
U1  Vout plot_v1		
U2  V1 plot_v1		
U3  V2 plot_v1		
v5  Z2 GND sine		
U4  Z2 plot_v1		
X1  Net-_R1-Pad2_ Vout Net-_X1-Pad3_ V1 GND Z2 GND GND V2 Net-_X1-Pad10_ MPY100		

.end
