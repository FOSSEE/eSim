* C:\eSim\eSim\src\SubcircuitLibrary\LOGIC_ADDER\LOGIC_ADDER.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/24/2018 7:23:20 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  A B Net-_U2-Pad3_ d_and		
U4  Net-_U3-Pad3_ CIN Net-_U4-Pad3_ d_and		
U3  A B Net-_U3-Pad3_ d_xor		
U5  Net-_U3-Pad3_ CIN SUM d_xor		
U6  Net-_U2-Pad3_ Net-_U4-Pad3_ CARRY d_or		
U1  A B CIN SUM CARRY PORT		

.end
