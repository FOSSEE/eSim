* D:\FOSSEE\eSim\library\SubcircuitLibrary\tff_1\tff_1.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/17/25 12:05:50

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ d_and		
U3  Net-_U1-Pad2_ Net-_U1-Pad1_ Net-_U3-Pad3_ d_and		
U4  Net-_U1-Pad3_ Net-_U2-Pad4_ Net-_U4-Pad3_ d_nand		
U5  Net-_U2-Pad5_ Net-_U3-Pad3_ Net-_U5-Pad3_ d_nand		
U6  Net-_U2-Pad6_ Net-_U4-Pad3_ Net-_U6-Pad3_ d_and		
U7  Net-_U5-Pad3_ Net-_U2-Pad3_ Net-_U7-Pad3_ d_and		
U8  Net-_U6-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ d_nand		
U9  Net-_U2-Pad5_ Net-_U7-Pad3_ Net-_U2-Pad4_ d_nand		
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ PORT		

.end
