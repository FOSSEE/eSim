.title KiCad schematic
R3 Net-_I1-Pad2_ Net-_Q3-Pad1_ 2k
Q6 Net-_Q4-Pad1_ Net-_I3-Pad1_ Net-_Q11-Pad2_ eSim_PNP
R2 Net-_Q4-Pad1_ Net-_I4-Pad1_ 50k
Q7 Net-_Q11-Pad2_ Net-_I4-Pad2_ Net-_Q3-Pad1_ eSim_NPN
R8 Net-_M4-Pad2_ Net-_I4-Pad1_ 10k
R7 Net-_M1-Pad2_ Net-_I4-Pad1_ 10k
R4 Net-_Q1-Pad1_ Net-_I4-Pad1_ 20k
Q8 Net-_Q1-Pad1_ Net-_I3-Pad1_ Net-_Q12-Pad2_ eSim_PNP
Q11 Net-_M1-Pad2_ Net-_Q11-Pad2_ Net-_I5-Pad1_ eSim_NPN
I4 Net-_I4-Pad1_ Net-_I4-Pad2_ 1m
I5 Net-_I5-Pad1_ Net-_I1-Pad2_ 500u
M2 Net-_M1-Pad1_ Net-_M1-Pad1_ Net-_I1-Pad2_ Net-_I1-Pad2_ eSim_MOS_N
M3 Net-_M3-Pad1_ Net-_M1-Pad1_ Net-_I1-Pad2_ Net-_I1-Pad2_ eSim_MOS_N
Q12 Net-_M4-Pad2_ Net-_Q12-Pad2_ Net-_I5-Pad1_ eSim_NPN
Q5 Net-_I3-Pad1_ Net-_I3-Pad1_ Net-_Q5-Pad3_ eSim_PNP
R1 Net-_Q5-Pad3_ Net-_I4-Pad1_ 50k
I1 Net-_Q1-Pad3_ Net-_I1-Pad2_ 400u
Q4 Net-_Q4-Pad1_ Net-_Q3-Pad2_ Net-_Q1-Pad3_ eSim_NPN
I3 Net-_I3-Pad1_ Net-_I1-Pad2_ 300u
I2 Net-_I4-Pad1_ Net-_Q2-Pad3_ 200u
U1 Net-_M3-Pad1_ Net-_I1-Pad2_ Net-_Q3-Pad2_ Net-_Q1-Pad2_ Net-_I4-Pad1_ PORT
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN
Q3 Net-_Q3-Pad1_ Net-_Q3-Pad2_ Net-_Q2-Pad3_ eSim_PNP
Q2 Net-_Q2-Pad1_ Net-_Q1-Pad2_ Net-_Q2-Pad3_ eSim_PNP
R5 Net-_I1-Pad2_ Net-_Q2-Pad1_ 2k
Q9 Net-_Q12-Pad2_ Net-_I4-Pad2_ Net-_Q2-Pad1_ eSim_NPN
R6 Net-_I1-Pad2_ Net-_Q10-Pad3_ 5k
Q10 Net-_I4-Pad2_ Net-_I4-Pad2_ Net-_Q10-Pad3_ eSim_NPN
M1 Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_I4-Pad1_ Net-_I4-Pad1_ eSim_MOS_P
M4 Net-_M3-Pad1_ Net-_M4-Pad2_ Net-_I4-Pad1_ Net-_I4-Pad1_ eSim_MOS_P
.end
