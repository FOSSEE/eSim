.title KiCad schematic
U4 Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ V_Y2 V_Y1 V_Y4 V_Y3 dac_bridge_4
U5 V_Y3 plot_v1
U6 V_Y4 plot_v1
v1 Net-_X1-Pad14_ GND 5
U7 Net-_V_B4-Pad1_ Net-_V_A4-Pad1_ Net-_V_B3-Pad1_ Net-_V_A3-Pad1_ Net-_U7-Pad5_ Net-_U7-Pad6_ Net-_U7-Pad7_ Net-_U7-Pad8_ adc_bridge_4
V_A1 Net-_V_A1-Pad1_ GND DC
V_A2 Net-_V_A2-Pad1_ GND DC
V_B1 Net-_V_B1-Pad1_ GND DC
V_B2 Net-_V_B2-Pad1_ GND DC
U2 Net-_V_A1-Pad1_ Net-_V_B1-Pad1_ Net-_V_A2-Pad1_ Net-_V_B2-Pad1_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ adc_bridge_4
V_A3 Net-_V_A3-Pad1_ GND DC
V_B3 Net-_V_B3-Pad1_ GND DC
V_B4 Net-_V_B4-Pad1_ GND DC
V_A4 Net-_V_A4-Pad1_ GND DC
X1 Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U4-Pad2_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U4-Pad1_ GND Net-_U4-Pad4_ Net-_U7-Pad8_ Net-_U7-Pad7_ Net-_U4-Pad3_ Net-_U7-Pad6_ Net-_U7-Pad5_ Net-_X1-Pad14_ 74HC00
U1 V_Y1 plot_v1
U3 V_Y2 plot_v1
.end
