* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Jun 22 15:31:09 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
X1  Net-_R2-Pad1_ In Out UA741		
R2  Net-_R2-Pad1_ GND 1k		
R3  GND Out 1k		
R5  Out In 1k		
v1  Net-_R1-Pad2_ GND sine		
R1  In Net-_R1-Pad2_ 1k		

.end
