.title KiCad schematic
R5 Net-_Q5-Pad3_ Net-_Q1-Pad3_ 1k
R3 Net-_Q1-Pad2_ Net-_Q1-Pad3_ 2k
Q6 Net-_Q5-Pad1_ Net-_Q4-Pad1_ Net-_Q6-Pad3_ eSim_NPN
Q5 Net-_Q5-Pad1_ Net-_Q5-Pad1_ Net-_Q5-Pad3_ eSim_PNP
U1 Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q10-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad1_ Net-_R6-Pad2_ Net-_R1-Pad1_ Net-_Q10-Pad3_ Net-_Q1-Pad3_ Net-_Q7-Pad1_ PORT
R7 Net-_Q7-Pad3_ Net-_Q1-Pad3_ 1k
Q9 Net-_Q1-Pad3_ Net-_Q7-Pad1_ Net-_Q10-Pad3_ eSim_NPN
Q7 Net-_Q7-Pad1_ Net-_Q5-Pad1_ Net-_Q7-Pad3_ eSim_PNP
D1 Net-_Q7-Pad1_ Net-_Q10-Pad2_ eSim_Diode
Q10 Net-_Q10-Pad1_ Net-_Q10-Pad2_ Net-_Q10-Pad3_ eSim_PNP
Q8 Net-_Q10-Pad2_ Net-_Q2-Pad1_ Net-_Q6-Pad3_ eSim_NPN
R6 Net-_Q10-Pad1_ Net-_R6-Pad2_ 1k
R2 Net-_Q2-Pad1_ Net-_Q10-Pad1_ 10k
R4 Net-_Q10-Pad1_ Net-_Q4-Pad1_ 10k
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_PNP
Q3 Net-_Q2-Pad3_ Net-_Q1-Pad1_ Net-_Q1-Pad2_ eSim_PNP
R1 Net-_R1-Pad1_ Net-_Q1-Pad1_ 200k
Q4 Net-_Q4-Pad1_ Net-_Q4-Pad2_ Net-_Q2-Pad3_ eSim_PNP
Q2 Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_PNP
.end
