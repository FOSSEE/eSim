* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/TC74HC4028AP/TC74HC4028AP.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Jul  5 21:40:54 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  /A_bar /B_bar /Gnd /Vd Net-_U1-Pad5_ /C_bar /D_bar Y0		
X4  /Vd /A /B_bar /Gnd /C_bar /D_bar Net-_U1-Pad10_ Y1		
X6  /Vd /A_bar /B /Gnd /C_bar /D_bar Net-_U1-Pad15_ Y2		
X9  /Vd /A /B /Gnd /C_bar /D_bar Net-_U1-Pad19_ Y3		
X2  /Vd /A_bar /B_bar /Gnd /C /D_bar Net-_U1-Pad7_ Y4		
X5  /Vd /A /B_bar /Gnd /C /D_bar Net-_U1-Pad13_ Y5		
X7  /Vd /A_bar /B /Gnd /C /D_bar Net-_U1-Pad16_ Y6		
X10  /Vd /A /B /Gnd /C /D_bar Net-_U1-Pad20_ Y7		
X8  /Vd /A /B_bar /Gnd /C_bar /D Net-_U1-Pad17_ Y9		
scmode1  SKY130mode		
U1  /Vd /A_bar /B_bar /D_bar Net-_U1-Pad5_ /A Net-_U1-Pad7_ /Gnd Net-_U1-Pad9_ Net-_U1-Pad10_ /C /C_bar Net-_U1-Pad13_ /B Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ /D Net-_U1-Pad19_ Net-_U1-Pad20_ PORT		
X3  /Vd /A_bar /B_bar /Gnd /C_bar /D Net-_U1-Pad9_ Y8		

.end
