* C:\Users\pavithra\eSim-Workspace\envelope_detector\envelope_detector.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/03/25 13:19:10

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_D1-Pad1_ GND sine		
D1  Net-_D1-Pad1_ Net-_C1-Pad1_ eSim_Diode		
C1  Net-_C1-Pad1_ GND 0.047u		
R1  Net-_C1-Pad1_ GND 10k		

.end
