* C:\FOSSEE\eSim\library\SubcircuitLibrary\SN55188\SN55188.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/09/25 00:32:09

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X2  Vcc+ Net-_U1-Pad2_ Net-_U1-Pad2_ gnd Vcc- Net-_U1-Pad3_ SN55188_0		
X3  Vcc+ Net-_U1-Pad9_ Net-_U1-Pad10_ gnd Vcc- Net-_U1-Pad8_ SN55188_0		
X1  Vcc+ Net-_U1-Pad4_ Net-_U1-Pad5_ gnd Vcc- Net-_U1-Pad6_ SN55188_0		
X4  Vcc+ Net-_U1-Pad12_ Net-_U1-Pad13_ gnd Vcc- Net-_U1-Pad11_ SN55188_0		
U1  Vcc- Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ gnd Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Vcc+ PORT		

.end
