* C:\Users\HP\eSim-Workspace\dualtimer\dualtimer.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/18/19 20:07:24

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R3-Pad2_ c1 Net-_C2-Pad1_ Net-_R1-Pad1_ out1 c1 GND c2 out2 Net-_R1-Pad1_ Net-_C3-Pad1_ c2 Net-_R5-Pad2_ Net-_R1-Pad1_ 556		
C2  Net-_C2-Pad1_ GND 0.001u		
C3  Net-_C3-Pad1_ GND 0.001u		
R4  Net-_R3-Pad2_ c1 100k		
R6  Net-_R5-Pad2_ c2 100k		
R3  Net-_R1-Pad1_ Net-_R3-Pad2_ 1k		
R5  Net-_R1-Pad1_ Net-_R5-Pad2_ 1k		
C1  c1 GND 100n		
C4  c2 GND 100n		
R1  Net-_R1-Pad1_ Net-_D1-Pad2_ 1000		
D1  out1 Net-_D1-Pad2_ LED		
R2  out1 Net-_D2-Pad2_ 1k		
D2  GND Net-_D2-Pad2_ LED		
R7  Net-_R1-Pad1_ Net-_D3-Pad2_ 1000		
D3  out2 Net-_D3-Pad2_ LED		
R8  out2 Net-_D4-Pad2_ 1k		
D4  GND Net-_D4-Pad2_ LED		
v1  Net-_R1-Pad1_ GND DC		
U3  c2 IC		
U2  c1 IC		
U4  out2 plot_v1		
U1  out1 plot_v1		
U6  c2 plot_v1		
U5  c1 plot_v1		

.end
