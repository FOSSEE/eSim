* /opt/eSim/src/SubcircuitLibrary/diac/diac.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Dec  8 15:35:49 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  1 2 PORT		
U1  1 1 2 aswitch		
U2  1 1 2 aswitch		

.end
