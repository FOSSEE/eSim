* C:\Users\Aditya\eSim-Workspace\SRAM\SRAM.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/24/24 12:32:19

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  WL GND pulse		
v2  BL GND pulse		
v3  Net-_X1-Pad1_ GND DC		
U1  WL plot_v1		
U2  BL plot_v1		
U5  NOT_BL plot_v1		
U4  Q plot_v1		
U3  NOT_Q plot_v1		
R1  NOT_Q GND 1000k		
R2  Q GND 1000k		
v4  NOT_BL GND pulse		
X1  Net-_X1-Pad1_ WL BL NOT_BL GND Q NOT_Q SRAM_Cell		

.end
