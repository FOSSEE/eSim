* C:\Users\senba\Desktop\FOSSEE\eSim\library\SubcircuitLibrary\SN74LS76\SN74LS76.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/10/25 06:29:32

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X2  Net-_U1-Pad6_ Net-_U3-Pad2_ Net-_U1-Pad5_ Net-_U2-Pad2_ 3_and		
X3  Net-_U1-Pad5_ Net-_U1-Pad4_ Net-_U1-Pad6_ Net-_U2-Pad1_ 3_and		
X4  Net-_U1-Pad1_ Net-_U4-Pad2_ Net-_U1-Pad2_ Net-_U5-Pad1_ 3_and		
X5  Net-_U1-Pad2_ Net-_U1-Pad4_ Net-_U1-Pad1_ Net-_U5-Pad2_ 3_and		
X1  Net-_U1-Pad5_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U3-Pad1_ 4_and		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ d_inverter		
X6  Net-_U1-Pad4_ Net-_U1-Pad7_ Net-_U1-Pad6_ Net-_U1-Pad1_ Net-_U4-Pad1_ 4_and		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ d_inverter		
U5  Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U1-Pad5_ d_nor		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad1_ d_nor		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ PORT		

.end
