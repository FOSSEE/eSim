* C:\FOSSEE\eSim\library\SubcircuitLibrary\SN74H55\SN74H55.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/21/25 12:33:56

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_X1-Pad5_ 4_and		
X2  Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ Net-_U3-Pad13_ Net-_X2-Pad5_ 4_and		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ d_inverter		
X3  Net-_X1-Pad5_ Net-_X2-Pad5_ Net-_U1-Pad2_ Net-_U3-Pad5_ Net-_U2-Pad1_ 4_OR		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ d_inverter		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U3-Pad5_ ? ? Net-_U2-Pad2_ Net-_U1-Pad1_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ Net-_U3-Pad13_ ? PORT		

.end
