* C:\Users\malli\eSim\src\SubcircuitLibrary\5_and\5_and.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/26/19 18:53:13

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U3-Pad1_ 3_and		
U2  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U2-Pad3_ d_and		
U3  Net-_U3-Pad1_ Net-_U2-Pad3_ Net-_U1-Pad6_ d_and		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ PORT		

.end
