* C:\FOSSEE\eSim\library\SubcircuitLibrary\SN55188_0\SN55188_0.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/05/25 19:31:16

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_D4-Pad2_ eSim_PNP		
Q2  Net-_Q1-Pad1_ Net-_Q2-Pad2_ Net-_D9-Pad1_ eSim_NPN		
Q3  Net-_D5-Pad1_ Net-_Q1-Pad1_ Net-_Q3-Pad3_ eSim_NPN		
Q5  Net-_D5-Pad2_ Net-_Q3-Pad3_ Net-_Q2-Pad2_ eSim_NPN		
R3  Net-_Q1-Pad1_ Net-_D9-Pad1_ 10k		
R1  Net-_D4-Pad2_ Net-_Q1-Pad2_ 3.6k		
D4  Net-_D3-Pad2_ Net-_D4-Pad2_ eSim_Diode		
D3  Net-_D1-Pad1_ Net-_D3-Pad2_ eSim_Diode		
R2  Net-_D8-Pad2_ Net-_D1-Pad1_ 8.2k		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
D2  Net-_D1-Pad1_ Net-_D2-Pad2_ eSim_Diode		
Q4  Net-_D8-Pad2_ Net-_D5-Pad1_ Net-_Q4-Pad3_ eSim_NPN		
R4  Net-_D8-Pad2_ Net-_D5-Pad1_ 6.2k		
R6  Net-_Q4-Pad3_ Net-_D6-Pad2_ 70		
D6  Net-_D5-Pad2_ Net-_D6-Pad2_ eSim_Diode		
D7  Net-_D6-Pad2_ Net-_D5-Pad2_ eSim_Diode		
D5  Net-_D5-Pad1_ Net-_D5-Pad2_ eSim_Diode		
R7  Net-_Q2-Pad2_ Net-_D9-Pad1_ 70		
R5  Net-_Q3-Pad3_ Net-_D9-Pad1_ 3.7k		
D9  Net-_D9-Pad1_ Net-_D6-Pad2_ eSim_Diode		
R8  Net-_D6-Pad2_ Net-_R8-Pad2_ 300		
D8  Net-_D6-Pad2_ Net-_D8-Pad2_ eSim_Diode		
U1  Net-_D8-Pad2_ Net-_D1-Pad2_ Net-_D2-Pad2_ Net-_Q1-Pad2_ Net-_D9-Pad1_ Net-_R8-Pad2_ PORT		

.end
