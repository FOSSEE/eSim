* C:\FOSSEE\eSim\library\SubcircuitLibrary\74HC27\74HC27.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/17/2025 4:51:11 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad2_ Net-_U1-Pad1_ Net-_U2-Pad3_ d_or		
U4  Net-_U2-Pad3_ Net-_U1-Pad3_ Net-_U4-Pad3_ d_or		
U6  Net-_U4-Pad3_ Net-_U1-Pad4_ d_inverter		
U13  Net-_U1-Pad12_ Net-_U1-Pad10_ Net-_U11-Pad1_ d_or		
U11  Net-_U11-Pad1_ Net-_U1-Pad8_ Net-_U11-Pad3_ d_or		
U9  Net-_U11-Pad3_ Net-_U1-Pad6_ d_inverter		
U12  Net-_U1-Pad11_ Net-_U1-Pad9_ Net-_U10-Pad1_ d_or		
U10  Net-_U10-Pad1_ Net-_U1-Pad7_ Net-_U10-Pad3_ d_or		
U8  Net-_U10-Pad3_ Net-_U1-Pad5_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ PORT		

.end
