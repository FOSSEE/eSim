* D:\FOSSEE\eSim\library\SubcircuitLibrary\TS391_IC\TS391_IC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/22/24 20:07:00

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
I1  Net-_I1-Pad1_ Net-_D2-Pad1_ 3.5u		
I2  Net-_I1-Pad1_ Net-_I2-Pad2_ 100u		
I3  Net-_I1-Pad1_ Net-_D3-Pad1_ 3.5u		
I4  Net-_I1-Pad1_ Net-_I4-Pad2_ 100u		
D2  Net-_D2-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q4  Net-_Q4-Pad1_ Net-_D3-Pad2_ Net-_I2-Pad2_ eSim_PNP		
Q2  Net-_Q2-Pad1_ Net-_D1-Pad2_ Net-_I2-Pad2_ eSim_PNP		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q1  Net-_Q1-Pad1_ Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_PNP		
Q3  Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_Q1-Pad1_ eSim_NPN		
Q5  Net-_Q4-Pad1_ Net-_Q2-Pad1_ Net-_Q1-Pad1_ eSim_NPN		
D3  Net-_D3-Pad1_ Net-_D3-Pad2_ eSim_Diode		
D4  Net-_D4-Pad1_ Net-_D3-Pad2_ eSim_Diode		
Q6  Net-_Q1-Pad1_ Net-_D4-Pad1_ Net-_D3-Pad2_ eSim_PNP		
Q7  Net-_I4-Pad2_ Net-_Q4-Pad1_ Net-_Q1-Pad1_ eSim_NPN		
Q8  Net-_Q8-Pad1_ Net-_I4-Pad2_ Net-_Q1-Pad1_ eSim_NPN		
R2  Net-_I1-Pad1_ Net-_Q8-Pad1_ 3.5k		
R1  Net-_R1-Pad1_ Net-_D4-Pad1_ 1k		
U1  Net-_Q8-Pad1_ Net-_Q1-Pad1_ Net-_R1-Pad1_ Net-_D1-Pad1_ Net-_I1-Pad1_ PORT		

.end
