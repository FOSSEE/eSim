* E:\FOSSEE\eSim\library\SubcircuitLibrary\SN54H87\SN54H87.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/02/25 08:58:06

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U10-Pad2_ d_inverter		
U3  Net-_U1-Pad2_ Net-_U3-Pad2_ d_inverter		
U11  Net-_U1-Pad3_ Net-_U10-Pad2_ Net-_U11-Pad3_ d_nand		
U4  Net-_U3-Pad2_ Net-_U13-Pad2_ d_inverter		
U9  Net-_U1-Pad4_ Net-_U10-Pad2_ Net-_U14-Pad1_ d_nand		
U7  Net-_U3-Pad2_ Net-_U14-Pad2_ d_inverter		
U10  Net-_U1-Pad5_ Net-_U10-Pad2_ Net-_U10-Pad3_ d_nand		
U8  Net-_U3-Pad2_ Net-_U15-Pad2_ d_inverter		
U5  Net-_U1-Pad6_ Net-_U10-Pad2_ Net-_U12-Pad1_ d_nand		
U6  Net-_U3-Pad2_ Net-_U12-Pad2_ d_inverter		
U13  Net-_U11-Pad3_ Net-_U13-Pad2_ Net-_U1-Pad10_ d_xor		
U14  Net-_U14-Pad1_ Net-_U14-Pad2_ Net-_U1-Pad9_ d_xor		
U15  Net-_U10-Pad3_ Net-_U15-Pad2_ Net-_U1-Pad7_ d_xor		
U12  Net-_U12-Pad1_ Net-_U12-Pad2_ Net-_U1-Pad8_ d_xor		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ GNDPWR GNDPWR GNDPWR GNDPWR PORT		

.end
