* C:\FOSSEE\eSim\library\SubcircuitLibrary\CD520b\CD520b.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/26/25 14:49:37

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U7  Net-_U7-Pad1_ Net-_U5-Pad3_ Net-_U1-Pad7_ Net-_U11-Pad4_ Net-_U7-Pad5_ Net-_U7-Pad1_ d_dff		
U9  Net-_U11-Pad2_ Net-_U7-Pad1_ Net-_U1-Pad7_ Net-_U11-Pad4_ Net-_U10-Pad1_ Net-_U11-Pad2_ d_dff		
U11  Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U1-Pad7_ Net-_U11-Pad4_ Net-_U11-Pad5_ Net-_U11-Pad1_ d_dff		
U13  Net-_U13-Pad1_ Net-_U11-Pad1_ Net-_U1-Pad7_ Net-_U11-Pad4_ Net-_U13-Pad5_ Net-_U13-Pad1_ d_dff		
U8  Net-_U7-Pad5_ Net-_U6-Pad1_ d_inverter		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ d_inverter		
U12  Net-_U11-Pad5_ Net-_U12-Pad2_ d_inverter		
U14  Net-_U13-Pad5_ Net-_U14-Pad2_ d_inverter		
U5  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U5-Pad3_ d_nand		
U6  Net-_U6-Pad1_ Net-_U10-Pad2_ Net-_U12-Pad2_ Net-_U14-Pad2_ Net-_U1-Pad5_ Net-_U1-Pad4_ Net-_U1-Pad3_ Net-_U1-Pad2_ dac_bridge_4		
U2  Net-_U1-Pad6_ Net-_U1-Pad8_ Net-_U2-Pad3_ Net-_U2-Pad4_ adc_bridge_2		
U3  Net-_U1-Pad1_ Net-_U3-Pad2_ adc_bridge_1		
U4  Net-_U3-Pad2_ Net-_U11-Pad4_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ PORT		

.end
