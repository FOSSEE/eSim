* C:\Users\Shanthipriya\Desktop\madeeasy\FOSSEE\eSim\library\SubcircuitLibrary\internal72\internal72.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/24/25 09:40:12

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U3-Pad1_ Net-_U1-Pad1_ Net-_U3-Pad3_ d_nand		
U4  Net-_U2-Pad2_ Net-_U4-Pad2_ Net-_U4-Pad3_ d_nand		
U5  Net-_U3-Pad3_ Net-_U4-Pad3_ Net-_U5-Pad3_ d_nand		
U2  Net-_U1-Pad3_ Net-_U2-Pad2_ d_inverter		
U7  Net-_U5-Pad3_ Net-_U1-Pad2_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U4-Pad2_ Net-_U3-Pad1_ d_dff		
U8  Net-_U4-Pad2_ Net-_U6-Pad2_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ d_dff		
U6  Net-_U1-Pad2_ Net-_U6-Pad2_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ ? ? Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ PORT		

.end
