* C:\Users\Shanthipriya\Desktop\madeeasy\FOSSEE\eSim\library\SubcircuitLibrary\f_origin\f_origin.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/10/25 01:12:40

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  /w /x /y /z Net-_U1-Pad5_ PORT		
U2  /y Net-_U2-Pad2_ d_inverter		
U3  /z Net-_U3-Pad2_ d_inverter		
X1  Net-_U4-Pad3_ Net-_U5-Pad3_ Net-_U6-Pad3_ Net-_U7-Pad3_ Net-_U1-Pad5_ 4_OR		
U4  Net-_U2-Pad2_ Net-_U3-Pad2_ Net-_U4-Pad3_ d_and		
U5  /x Net-_U2-Pad2_ Net-_U5-Pad3_ d_and		
U6  /x Net-_U3-Pad2_ Net-_U6-Pad3_ d_and		
U7  /w Net-_U2-Pad2_ Net-_U7-Pad3_ d_and		

.end
