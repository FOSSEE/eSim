* C:\Users\Shanthipriya\eSim-Workspace\7447\7447.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/11/25 02:00:36

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  W GND pulse		
v2  X GND pulse		
v3  Y GND pulse		
v4  Z GND pulse		
v5  Net-_X1-Pad5_ GND DC		
v6  Net-_X1-Pad6_ GND DC		
v7  Net-_X1-Pad7_ GND DC		
U1  Z plot_v1		
U2  Y plot_v1		
U3  X plot_v1		
U4  W plot_v1		
U5  a plot_v1		
U6  b plot_v1		
U7  c plot_v1		
U8  d plot_v1		
U9  e plot_v1		
U10  f plot_v1		
U11  g plot_v1		
X1  W X Y Z Net-_X1-Pad5_ Net-_X1-Pad6_ Net-_X1-Pad7_ a b c d e f g ? ? 74_48		

.end
