* C:\FOSSEE\eSim\library\SubcircuitLibrary\LOG_Amplifier\LOG_Amplifier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 9/11/2022 7:52:59 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  ? /Inp1 GND /Vneg ? Net-_Q1-Pad3_ /Vpos ? lm_741		
X2  ? /Inp2 GND /Vneg ? /Vout /Vpos ? lm_741		
Q1  /Inp1 Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
Q2  /Inp2 GND Net-_Q1-Pad3_ eSim_NPN		
R1  /Vout Net-_Q1-Pad2_ 3.2k		
R2  Net-_Q1-Pad2_ GND 5k		
C1  /Vout /Inp2 3.4u		
U1  /Inp1 /NC /Vout /Vpos /Vneg GND /NC /Inp2 PORT		

.end
