* eeschema netlist version 1.1 (spice format) creation date: wednesday 29 april 2015 05:48:14 pm ist
.include mos_n.lib
.include mos_p.lib

v1 in gnd  dc 5
m2 out in gnd gnd mos_n M=100u L=100u W=100u
m1 out in vcc vcc mos_p M=100u L=100u W=100u
c1  out gnd 1u
v2 vcc gnd  dc 5
* Plotting option vplot8_1

.tran  10e-03 100e-03 0e-03
.plot v(in) v(out) 
.end
