* /home/fossee/UpdatedExamples/HalfwaveRectifier_SCR/HalfwaveRectifier_SCR.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Mar  3 22:33:43 2016

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  in GND sine		
v2  pulse GND pulse		
R1  in A 100		
U2  in A plot_v2		
U1  in plot_v1		
U3  pulse plot_v1		
X1  GND pulse A SCR		

.end
