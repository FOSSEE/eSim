* eeschema netlist version 1.1 (spice format) creation date: 10/08/14 11:31:43
.include scr.sub

v2  2 0 pulse(0 5 4m 0 0 1m 20m)
* Plotting option vplot1
* Plotting option vplot
x3  0 2 4 scr
r1  4 1 500
v1  1 0 sine(0 100 50 0 0)

.tran  20e-06 20e-03 0e-00
.plot v(1)
.plot v(1)-v(4)
.end
