* C:\FOSSEE\eSim\library\SubcircuitLibrary\HD74HC30\HD74HC30.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/09/25 15:20:42

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U2-Pad1_ 4_and		
X2  Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U2-Pad2_ 4_and		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ d_and		
U3  Net-_U2-Pad3_ Net-_U1-Pad8_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ ? Net-_U1-Pad8_ ? ? Net-_U1-Pad11_ Net-_U1-Pad12_ ? ? PORT		

.end
