* C:\Users\Shanthipriya\eSim-Workspace\4_bit_FA\4_bit_FA.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/08/25 10:08:09

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  C0 plot_v1		
U3  A1 plot_v1		
U4  A2 plot_v1		
U5  A3 plot_v1		
U7  A4 plot_v1		
U1  B1 plot_v1		
U6  B4 plot_v1		
U8  B3 plot_v1		
U9  B2 plot_v1		
U10  S1 plot_v1		
U11  S2 plot_v1		
U12  S3 plot_v1		
U13  S4 plot_v1		
U14  C_out plot_v1		
X1  A1 B1 C0 A2 B2 A3 B3 A4 B4 S1 S2 S3 S4 C_out ? ? 283		
v1  C0 GND pulse		
v2  A1 GND pulse		
v3  A2 GND pulse		
v4  A3 GND pulse		
v5  A4 GND pulse		
v6  B1 GND pulse		
v7  B2 GND pulse		
v8  B3 GND pulse		
v9  B4 GND pulse		

.end
