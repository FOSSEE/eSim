* C:\FOSSEE\eSim\library\SubcircuitLibrary\SN74H62\SN74H62.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/10/25 11:11:56

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ d_and		
X1  Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U3-Pad5_ Net-_X1-Pad4_ 3_and		
X2  Net-_U3-Pad9_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_X2-Pad4_ 3_and		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ d_and		
X3  Net-_U1-Pad3_ Net-_X1-Pad4_ Net-_X2-Pad4_ Net-_U2-Pad3_ Net-_U3-Pad8_ 4_OR		
U4  Net-_U3-Pad8_ Net-_U3-Pad6_ d_inverter		
U3  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U3-Pad5_ Net-_U3-Pad6_ ? Net-_U3-Pad8_ Net-_U3-Pad9_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U2-Pad1_ Net-_U2-Pad2_ ? PORT		

.end
