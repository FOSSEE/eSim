* D:\FOSSEE\eSim\library\SubcircuitLibrary\ref5010_2\ref5010_2.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/09/25 17:52:34

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  ? Net-_R1-Pad2_ Net-_R3-Pad2_ Net-_X1-Pad4_ ? Net-_R2-Pad2_ Net-_X1-Pad7_ ? lm_741		
R2  Net-_R1-Pad2_ Net-_R2-Pad2_ 1k		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 1k		
R3  Net-_R3-Pad1_ Net-_R3-Pad2_ 10k		
R4  Net-_R3-Pad2_ Net-_R4-Pad2_ 1k		
U1  Net-_I1-Pad2_ ? Net-_R2-Pad2_ ? ? Net-_R4-Pad2_ Net-_I1-Pad1_ Net-_R1-Pad1_ PORT		
v1  Net-_R3-Pad1_ Net-_R1-Pad1_ 1.2v		
I1  Net-_I1-Pad1_ Net-_I1-Pad2_ 0.000001		
R5  Net-_I1-Pad1_ Net-_R1-Pad1_ 60k		
v2  Net-_X1-Pad7_ GND 12v		
v3  Net-_X1-Pad4_ GND 12v		

.end
