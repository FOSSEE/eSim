* C:\esim\eSim\src\SubcircuitLibrary\5bit-Ripple_carry_adder\5bit-Ripple_carry_adder.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/23/19 02:16:47

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X4  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_X4-Pad3_ Net-_U1-Pad4_ ? Full-Adder		
X5  Net-_U1-Pad3_ Net-_U1-Pad5_ Net-_X5-Pad3_ Net-_U1-Pad7_ Net-_X4-Pad3_ Full-Adder		
X6  Net-_U1-Pad6_ Net-_U1-Pad8_ Net-_X6-Pad3_ Net-_U1-Pad10_ Net-_X5-Pad3_ Full-Adder		
X7  Net-_U1-Pad9_ Net-_U1-Pad11_ Net-_X7-Pad3_ Net-_U1-Pad13_ Net-_X6-Pad3_ Full-Adder		
X8  Net-_U1-Pad12_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_X7-Pad3_ Full-Adder		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ PORT		

.end
