* C:\Users\Shanthipriya\eSim-Workspace\13_nand_ic5\13_nand_ic5.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/29/25 16:11:34

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U9  A1 A2 A3 A4 A5 A6 A7 A8 Net-_U9-Pad9_ Net-_U9-Pad10_ Net-_U9-Pad11_ Net-_U9-Pad12_ Net-_U9-Pad13_ Net-_U9-Pad14_ Net-_U9-Pad15_ Net-_U9-Pad16_ adc_bridge_8		
U13  Net-_U13-Pad1_ OUT dac_bridge_1		
v1  A1 GND pulse		
v2  A2 GND pulse		
v3  A3 GND pulse		
v4  A4 GND pulse		
v5  A5 GND pulse		
v6  A6 GND pulse		
v7  A7 GND pulse		
v8  A8 GND pulse		
U17  OUT plot_v1		
U1  A1 plot_v1		
U2  A2 plot_v1		
U3  A3 plot_v1		
U4  A4 plot_v1		
U5  A5 plot_v1		
U6  A6 plot_v1		
U7  A7 plot_v1		
U8  A8 plot_v1		
U10  A9 A10 A11 A12 A13 Net-_U10-Pad6_ Net-_U10-Pad7_ Net-_U10-Pad8_ Net-_U10-Pad9_ Net-_U10-Pad10_ adc_bridge_5		
v9  A9 GND pulse		
v10  A10 GND pulse		
v11  A11 GND pulse		
v12  A12 GND pulse		
v13  A13 GND pulse		
U11  A13 plot_v1		
U12  A12 plot_v1		
U14  A11 plot_v1		
U15  A10 plot_v1		
U16  A9 plot_v1		
X1  Net-_U9-Pad9_ Net-_U9-Pad10_ Net-_U9-Pad11_ Net-_U9-Pad12_ Net-_U9-Pad13_ Net-_U9-Pad14_ Net-_U9-Pad15_ Net-_U9-Pad16_ Net-_U10-Pad6_ Net-_U10-Pad7_ Net-_U10-Pad8_ Net-_U10-Pad9_ Net-_U10-Pad10_ Net-_U13-Pad1_ 133		

.end
