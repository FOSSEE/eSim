* C:\FOSSEE\eSim\library\SubcircuitLibrary\CD4069\CD4069.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/04/22 15:25:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M9  Net-_M10-Pad1_ Net-_M10-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_P		
M10  Net-_M10-Pad1_ Net-_M10-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad3_ eSim_MOS_N		
M11  Net-_M11-Pad1_ Net-_M11-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_P		
M12  Net-_M11-Pad1_ Net-_M11-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad3_ eSim_MOS_N		
M5  Net-_M5-Pad1_ Net-_M5-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_P		
M6  Net-_M5-Pad1_ Net-_M5-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad3_ eSim_MOS_N		
M7  Net-_M7-Pad1_ Net-_M7-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_P		
M8  Net-_M7-Pad1_ Net-_M7-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad3_ eSim_MOS_N		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_P		
M2  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad3_ eSim_MOS_N		
M3  Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_P		
M4  Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M10-Pad3_ Net-_M10-Pad3_ eSim_MOS_N		
U1  Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M5-Pad2_ Net-_M5-Pad1_ Net-_M10-Pad2_ Net-_M10-Pad1_ Net-_M10-Pad3_ Net-_M11-Pad1_ Net-_M11-Pad2_ Net-_M7-Pad1_ Net-_M7-Pad2_ Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ PORT		

.end
