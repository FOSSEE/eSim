* C:\FOSSEE\eSim\library\SubcircuitLibrary\lm3909\lm3909.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/09/25 19:06:02

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
R1  Net-_R1-Pad1_ Net-_Q1-Pad1_ 12		
R4  Net-_D1-Pad1_ Net-_Q1-Pad3_ 20k		
R2  Net-_R2-Pad1_ Net-_R2-Pad2_ 6k		
R3  Net-_R2-Pad2_ Net-_D1-Pad1_ 3k		
R5  Net-_Q1-Pad2_ Net-_Q2-Pad2_ 20k		
R6  Net-_Q2-Pad2_ Net-_Q1-Pad3_ 10k		
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
R7  Net-_Q2-Pad3_ Net-_R2-Pad1_ 100		
R8  Net-_Q1-Pad1_ Net-_Q1-Pad2_ 400		
R9  Net-_Q1-Pad2_ Net-_D1-Pad2_ 400		
Q3  Net-_D1-Pad2_ Net-_Q3-Pad2_ Net-_D1-Pad1_ eSim_NPN		
U1  Net-_R2-Pad2_ Net-_D1-Pad2_ ? Net-_D1-Pad1_ Net-_Q1-Pad1_ Net-_R1-Pad1_ ? Net-_R2-Pad1_ PORT		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q5  Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_Q1-Pad1_ eSim_PNP		
Q4  Net-_Q3-Pad2_ Net-_Q2-Pad1_ Net-_Q1-Pad1_ eSim_PNP		

.end
