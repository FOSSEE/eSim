* C:\eSim\eSim\src\SubcircuitLibrary\MUX\MUX.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/24/2018 7:29:10 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U1-Pad2_ Net-_U2-Pad2_ Net-_U3-Pad3_ d_and		
U4  Net-_U1-Pad1_ Net-_U1-Pad3_ Net-_U4-Pad3_ d_and		
U5  Net-_U3-Pad3_ Net-_U4-Pad3_ Net-_U1-Pad4_ d_or		
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ PORT		

.end
