.title KiCad schematic
U1 Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad11_ PORT
U19 Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U19-Pad3_ d_and
U20 Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U20-Pad3_ d_and
U23 Net-_U21-Pad3_ Net-_U1-Pad11_ d_inverter
U21 Net-_U17-Pad3_ Net-_U18-Pad3_ Net-_U21-Pad3_ d_and
U24 Net-_U22-Pad3_ Net-_U1-Pad9_ d_inverter
U22 Net-_U19-Pad3_ Net-_U20-Pad3_ Net-_U22-Pad3_ d_and
U18 Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U18-Pad3_ d_and
U17 Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U17-Pad3_ d_and
.end
