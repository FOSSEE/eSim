* D:\FOSSEE\eSim\library\SubcircuitLibrary\TL331\TL331.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/12/24 00:57:13

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
D2  Net-_D2-Pad1_ Net-_D1-Pad2_ 10u		
I2  Net-_I1-Pad1_ Net-_I2-Pad2_ 80u		
D3  Net-_D3-Pad1_ Net-_D3-Pad2_ 10u		
Q2  Net-_Q2-Pad1_ Net-_D1-Pad2_ Net-_I2-Pad2_ eSim_PNP		
Q5  Net-_Q4-Pad1_ Net-_D3-Pad2_ Net-_I2-Pad2_ eSim_PNP		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q1  GND Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_PNP		
D4  Net-_D4-Pad1_ Net-_D3-Pad2_ eSim_Diode		
Q6  GND Net-_D4-Pad1_ Net-_D3-Pad2_ eSim_PNP		
I4  Net-_I1-Pad1_ Net-_I4-Pad2_ 80u		
Q3  Net-_Q2-Pad1_ Net-_Q2-Pad1_ Net-_Q3-Pad3_ eSim_NPN		
Q4  Net-_Q4-Pad1_ Net-_Q2-Pad1_ Net-_Q3-Pad3_ eSim_NPN		
Q7  Net-_I4-Pad2_ Net-_Q4-Pad1_ Net-_Q3-Pad3_ eSim_NPN		
Q8  Net-_Q8-Pad1_ Net-_I4-Pad2_ Net-_Q3-Pad3_ eSim_NPN		
R1  Net-_I1-Pad1_ Net-_Q8-Pad1_ 300		
I1  Net-_I1-Pad1_ Net-_D2-Pad1_ 80u		
I3  Net-_I1-Pad1_ Net-_D3-Pad1_ 80u		
U1  Net-_D1-Pad1_ Net-_D4-Pad1_ Net-_Q3-Pad3_ Net-_I1-Pad1_ Net-_Q8-Pad1_ PORT		

.end
