* C:\Users\senba\eSim-Workspace\74HC279_test\74HC279_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 12/17/25 11:39:14

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U3-Pad5_ Net-_U3-Pad6_ Net-_U3-Pad7_ Net-_U3-Pad5_ Net-_U3-Pad8_ Net-_U4-Pad1_ Net-_U4-Pad2_ 74HC279		
U3  Rbar Sbar Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U3-Pad5_ Net-_U3-Pad6_ Net-_U3-Pad7_ Net-_U3-Pad8_ adc_bridge_4		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Q Q1 dac_bridge_2		
v1  Rbar GND pulse		
v2  Sbar GND pulse		
v3  Net-_U3-Pad3_ GND pulse		
v4  Net-_U3-Pad4_ GND pulse		
U5  Q plot_v1		
U6  Q1 plot_v1		
U1  Rbar plot_v1		
U2  Sbar plot_v1		

.end
