* C:\Users\Chaithu\FOSSEE\eSim\library\SubcircuitLibrary\sn54als29827\sn54als29827.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 5/28/2025 9:43:02 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U10-Pad2_ d_and		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U1-Pad18_ Net-_U1-Pad19_ Net-_U1-Pad20_ Net-_U1-Pad21_ Net-_U1-Pad22_ PORT		
U3  Net-_U1-Pad4_ Net-_U10-Pad2_ Net-_U1-Pad14_ tristate_buff		
U5  Net-_U1-Pad3_ Net-_U10-Pad2_ Net-_U1-Pad13_ tristate_buff		
U4  Net-_U1-Pad6_ Net-_U10-Pad2_ Net-_U1-Pad16_ tristate_buff		
U6  Net-_U1-Pad7_ Net-_U10-Pad2_ Net-_U1-Pad22_ tristate_buff		
U7  Net-_U1-Pad10_ Net-_U10-Pad2_ Net-_U1-Pad17_ tristate_buff		
U8  Net-_U1-Pad8_ Net-_U10-Pad2_ Net-_U1-Pad15_ tristate_buff		
U9  Net-_U1-Pad5_ Net-_U10-Pad2_ Net-_U1-Pad18_ tristate_buff		
U10  Net-_U1-Pad9_ Net-_U10-Pad2_ Net-_U1-Pad19_ tristate_buff		
U11  Net-_U1-Pad11_ Net-_U10-Pad2_ Net-_U1-Pad21_ tristate_buff		
U12  Net-_U1-Pad12_ Net-_U10-Pad2_ Net-_U1-Pad20_ tristate_buff		

.end
