* /home/kamalesh/Downloads/eSim-2.3/library/SubcircuitLibrary/oscillator_driver/oscillator_driver.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Apr  5 18:48:44 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_C101-Pad2_ Net-_C101-Pad2_ mosfet_n		
M2  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M3  Net-_M3-Pad1_ Net-_M1-Pad1_ Net-_C101-Pad2_ Net-_C101-Pad2_ mosfet_n		
M4  Net-_M3-Pad1_ Net-_M1-Pad1_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M5  Net-_M5-Pad1_ Net-_M3-Pad1_ Net-_C101-Pad2_ Net-_C101-Pad2_ mosfet_n		
M6  Net-_M5-Pad1_ Net-_M3-Pad1_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
M7  Net-_C101-Pad1_ Net-_M5-Pad1_ Net-_C101-Pad2_ Net-_C101-Pad2_ mosfet_n		
M8  Net-_C101-Pad1_ Net-_M5-Pad1_ Net-_M2-Pad3_ Net-_M2-Pad3_ mosfet_p		
U1  ? Net-_C101-Pad2_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M2-Pad3_ Net-_C101-Pad1_ PORT		
C101  Net-_C101-Pad1_ Net-_C101-Pad2_ 1u		

.end
