.title KiCad schematic
U1 Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ GND Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ GND Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT
X2 Net-_U1-Pad12_ Net-_U5-Pad2_ Net-_U1-Pad2_ Net-_U7-Pad1_ 3_and
X3 Net-_U1-Pad12_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U7-Pad2_ 3_and
U7 Net-_U7-Pad1_ Net-_U7-Pad2_ Net-_U1-Pad13_ d_nor
X4 Net-_U1-Pad1_ Net-_U1-Pad14_ Net-_U1-Pad13_ Net-_U1-Pad2_ Net-_U6-Pad1_ 4_and
U6 Net-_U6-Pad1_ Net-_U3-Pad1_ d_inverter
U12 Net-_U12-Pad1_ Net-_U12-Pad2_ d_inverter
X7 Net-_U1-Pad9_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U13-Pad2_ 3_and
X6 Net-_U1-Pad9_ Net-_U11-Pad2_ Net-_U1-Pad6_ Net-_U13-Pad1_ 3_and
X1 Net-_U1-Pad12_ Net-_U1-Pad3_ Net-_U1-Pad1_ Net-_U5-Pad1_ 3_and
U5 Net-_U5-Pad1_ Net-_U5-Pad2_ d_inverter
U3 Net-_U3-Pad1_ Net-_U1-Pad13_ Net-_U2-Pad2_ d_and
U2 Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U1-Pad12_ d_nor
U4 Net-_U1-Pad1_ Net-_U1-Pad13_ Net-_U2-Pad1_ d_and
U9 Net-_U12-Pad2_ Net-_U1-Pad8_ Net-_U8-Pad2_ d_and
U8 Net-_U10-Pad3_ Net-_U8-Pad2_ Net-_U1-Pad9_ d_nor
U11 Net-_U11-Pad1_ Net-_U11-Pad2_ d_inverter
X5 Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad5_ Net-_U11-Pad1_ 3_and
U10 Net-_U1-Pad5_ Net-_U1-Pad8_ Net-_U10-Pad3_ d_and
U13 Net-_U13-Pad1_ Net-_U13-Pad2_ Net-_U1-Pad8_ d_nor
X8 Net-_U1-Pad5_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad6_ Net-_U12-Pad1_ 4_and
.end
