.title KiCad schematic
R8 Net-_D4-Pad1_ Net-_D5-Pad2_ 1k
R4 Net-_Q5-Pad2_ Net-_D5-Pad2_ 4k
R5 Net-_D2-Pad2_ Net-_D5-Pad2_ 2.5k
Q7 Net-_Q7-Pad1_ Net-_D2-Pad2_ Net-_D2-Pad2_ eSim_NPN
D4 Net-_D4-Pad1_ Net-_D2-Pad2_ eSim_Diode
R7 GND Net-_Q12-Pad2_ 625
Q12 Net-_D5-Pad1_ Net-_Q12-Pad2_ GND eSim_NPN
Q9 Net-_D4-Pad1_ Net-_Q7-Pad1_ Net-_Q12-Pad2_ eSim_NPN
Q4 Net-_D2-Pad2_ Net-_Q2-Pad3_ GND eSim_NPN
R3 GND Net-_Q2-Pad3_ 1.6k
D1 GND Net-_D1-Pad2_ eSim_Diode
U1 Net-_D1-Pad2_ Net-_D2-Pad2_ Net-_D5-Pad1_ PORT
D6 Net-_D6-Pad1_ GND eSim_Diode
D2 Net-_D2-Pad1_ Net-_D2-Pad2_ eSim_Diode
Q2 Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_NPN
Q3 Net-_D5-Pad2_ Net-_Q2-Pad1_ Net-_D2-Pad1_ eSim_NPN
Q13 Net-_Q2-Pad2_ Net-_Q1-Pad1_ Net-_D6-Pad1_ eSim_NPN
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_D1-Pad2_ eSim_NPN
R1 Net-_Q1-Pad2_ Net-_D5-Pad2_ 4k
R2 Net-_Q2-Pad1_ Net-_D5-Pad2_ 2.5k
R11 Net-_Q2-Pad2_ Net-_D5-Pad2_ 4.25k
v1 Net-_D5-Pad2_ GND 5
R10 Net-_Q10-Pad1_ Net-_D5-Pad2_ 85
Q11 Net-_Q10-Pad1_ Net-_Q10-Pad3_ Net-_D5-Pad1_ eSim_NPN
D5 Net-_D5-Pad1_ Net-_D5-Pad2_ eSim_Diode
R9 Net-_Q12-Pad2_ Net-_Q10-Pad3_ 4k
Q10 Net-_Q10-Pad1_ Net-_D4-Pad1_ Net-_Q10-Pad3_ eSim_NPN
Q6 Net-_D2-Pad2_ Net-_Q5-Pad1_ Net-_Q6-Pad3_ eSim_NPN
R6 GND Net-_Q6-Pad3_ 1.6k
D3 GND Net-_D2-Pad2_ eSim_Diode
Q5 Net-_Q5-Pad1_ Net-_Q5-Pad2_ Net-_D2-Pad2_ eSim_NPN
Q8 Net-_Q7-Pad1_ Net-_Q6-Pad3_ GND eSim_NPN
.end
