* C:\FOSSEE\eSim\library\SubcircuitLibrary\SRAM_Cell\SRAM_Cell.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/27/24 10:55:15

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M1-Pad3_ Net-_M2-Pad2_ Net-_M1-Pad4_ Net-_M1-Pad4_ mosfet_n		
M4  Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad4_ Net-_M1-Pad4_ mosfet_n		
M6  Net-_M6-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad2_ Net-_M1-Pad4_ mosfet_n		
M2  Net-_M2-Pad1_ Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M2-Pad1_ mosfet_p		
M5  Net-_M2-Pad1_ Net-_M1-Pad3_ Net-_M2-Pad2_ Net-_M2-Pad1_ mosfet_p		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad4_ mosfet_n		
U1  Net-_M2-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M6-Pad1_ Net-_M1-Pad4_ Net-_M1-Pad3_ Net-_M2-Pad2_ PORT		

.end
