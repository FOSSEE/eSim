.title KiCad schematic
U1 Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ GND Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ GND PORT
U15 Net-_U12-Pad3_ Net-_U1-Pad13_ d_inverter
U17 Net-_U13-Pad3_ Net-_U1-Pad10_ d_inverter
U13 Net-_U13-Pad1_ Net-_U13-Pad2_ Net-_U13-Pad3_ d_nand
U9 Net-_U1-Pad9_ Net-_U13-Pad2_ d_inverter
U3 Net-_U1-Pad12_ Net-_U12-Pad2_ d_inverter
U12 Net-_U12-Pad1_ Net-_U12-Pad2_ Net-_U12-Pad3_ d_nand
U2 Net-_U1-Pad11_ Net-_U12-Pad1_ d_inverter
U8 Net-_U1-Pad8_ Net-_U13-Pad1_ d_inverter
U5 Net-_U1-Pad6_ Net-_U11-Pad2_ d_inverter
U7 Net-_U1-Pad5_ Net-_U11-Pad1_ d_inverter
U11 Net-_U11-Pad1_ Net-_U11-Pad2_ Net-_U11-Pad3_ d_nand
U10 Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ d_nand
U14 Net-_U11-Pad3_ Net-_U1-Pad4_ d_inverter
U16 Net-_U10-Pad3_ Net-_U1-Pad1_ d_inverter
U4 Net-_U1-Pad3_ Net-_U10-Pad2_ d_inverter
U6 Net-_U1-Pad2_ Net-_U10-Pad1_ d_inverter
.end
