* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/NAND_Latch/NAND_Latch.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sat Jun 14 10:44:18 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_X1-Pad4_ CMOS_INVTR		
X2  Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_X2-Pad4_ CMOS_INVTR		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ PORT		
X3  Net-_X1-Pad4_ Net-_U1-Pad4_ Net-_U1-Pad3_ Net-_U1-Pad5_ Net-_X3-Pad5_ NOR_2		
X4  Net-_X2-Pad4_ Net-_U1-Pad4_ Net-_U1-Pad3_ Net-_X3-Pad5_ Net-_U1-Pad5_ NOR_2		
scmode1  SKY130mode		

.end
