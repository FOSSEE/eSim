* C:\FOSSEE\eSim\library\SubcircuitLibrary\MC14016B\MC14016B.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/23/25 15:06:49

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ d_inverter		
U2  Net-_U1-Pad2_ Net-_U2-Pad2_ d_inverter		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad4_ eSim_MOS_P		
M2  Net-_M1-Pad1_ Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M2-Pad4_ eSim_MOS_N		
U3  Net-_U2-Pad2_ Net-_M1-Pad2_ dac_bridge_1		
U5  Net-_M1-Pad3_ Net-_U1-Pad1_ Net-_M1-Pad1_ Net-_M1-Pad4_ Net-_M2-Pad4_ PORT		
U4  Net-_U1-Pad2_ Net-_M2-Pad2_ dac_bridge_1		

.end
