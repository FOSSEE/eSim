* /home/fossee/UpdatedExamples/Parallel_Resonance/Parallel_Resonance.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Mar  3 22:48:00 2016

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  out GND 100		
L1  out GND 100m		
C1  GND out 10u		
v1  in GND AC		
R2  out in 1000		
U1  in plot_v1		
U3  out plot_v1		

.end
