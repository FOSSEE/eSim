* eeschema netlist version 1.1 (spice format) creation date: 09/08/14 10:24:20
.include diode.lib
.include scr.sub

v1  1 2 sine(0 200 100 0 0)
v2  4 0 pulse(0 5 2m 0 0 1m 5m)
r1  5 3 500
x1  0 4 5 scr
d4  0 2 diode
d3  2 3 diode
d2  0 1 diode
d1  1 3 diode

.tran  10e-06 20e-03 0e-00
.plot v(1)-v(2) v(3)-v(5) 
.end
