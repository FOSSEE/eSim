* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/or_2/or_2.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Jul 10 18:26:57 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ PORT		
scmode1  SKY130mode		
X1  Net-_U1-Pad1_ Net-_U1-Pad4_ Net-_U1-Pad3_ Net-_U1-Pad2_ Net-_X1-Pad5_ NOR_2		
X2  Net-_X1-Pad5_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ CMOS_INVTR		

.end
