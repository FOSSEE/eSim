*** XSPICE_PWM for audio demo *****************************
* sin in --> pwm --> filter --> sin out to load

* PWM with input frequency 1200k, variable duty cycle
apwm in dout pwm
.model pwm d_pwm(
+ frequency = 1.2Meg
+ cntl_array = [-1 -0.99 0.99 1]
+ dc_array = [0.01 0.01 0.99 0.99]
+ init_phase = 90)

* D to A including inverted output
aout [~dout dout] [outn outp] dac1

.model dac1 dac_bridge(out_low = 0 out_high = 1 out_undef = 0
+ input_load = 5.0e-12 t_rise = 2e-9
+ t_fall = 2e-9)

* LC filter *********************
L1 outn outflcn 33u
CLfiltern outflcn 0 0.1u

Cboth outflcn outflcp 0.47u

L2 outp outflcp 33u
CLfilterp outflcp 0 0.1u
*********************************

* load
RLooad  outflcp  outflcn 8

* input voltage
Vin in 0 dc 0 sin (0 0.95 1.01k)
* reference for comparison (input shifted by 3.05 degrees for compensating latency)
Vref ref 0 dc 0 sin (0 0.95 1.01k 0 0 -3.05)

.control
tran 0.5u 20m uic
rusage
plot v(outn) v(outp) v(in)+2 xlimit 11.65m 12.15m ylabel 'digital output versus vin'
plot 0.99 * v(ref) - v(outflcp) + v(outflcn) ylimit -2m 2m ylabel 'Difference between input and output'
plot 0.99 * v(ref) v(outflcp)-v(outflcn)  ylabel 'Input and output'
.endc

.end
