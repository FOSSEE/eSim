* C:\Users\malli\eSim\src\SubcircuitLibrary\AD620\AD620.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/04/19 16:16:13

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X2  Net-_R8-Pad1_ Net-_R1-Pad2_ Net-_U1-Pad2_ Net-_R10-Pad2_ Net-_R10-Pad1_ Net-_R1-Pad1_ Net-_U1-Pad7_ ? lm_741		
X1  Net-_R7-Pad2_ Net-_R2-Pad1_ Net-_U1-Pad3_ Net-_R10-Pad2_ Net-_R9-Pad2_ Net-_R2-Pad2_ Net-_U1-Pad7_ ? lm_741		
X3  Net-_R11-Pad2_ Net-_R4-Pad1_ Net-_R3-Pad1_ Net-_R10-Pad2_ Net-_R12-Pad2_ Net-_R6-Pad1_ Net-_U1-Pad7_ ? lm_741		
R1  Net-_R1-Pad1_ Net-_R1-Pad2_ 24.7k		
R2  Net-_R2-Pad1_ Net-_R2-Pad2_ 24.7k		
R4  Net-_R4-Pad1_ Net-_R1-Pad1_ 10k		
R3  Net-_R3-Pad1_ Net-_R2-Pad2_ 10k		
R6  Net-_R6-Pad1_ Net-_R4-Pad1_ 10k		
R5  Net-_R5-Pad1_ Net-_R3-Pad1_ 10k		
U1  Net-_R1-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_R10-Pad2_ Net-_R5-Pad1_ Net-_R6-Pad1_ Net-_U1-Pad7_ Net-_R2-Pad1_ PORT		
R8  Net-_R8-Pad1_ Net-_R10-Pad2_ 0.297k		
R10  Net-_R10-Pad1_ Net-_R10-Pad2_ 1k		
R7  Net-_R10-Pad2_ Net-_R7-Pad2_ 0.297k		
R9  Net-_R10-Pad2_ Net-_R9-Pad2_ 1k		
R12  Net-_R10-Pad2_ Net-_R12-Pad2_ 1k		
R11  Net-_R10-Pad2_ Net-_R11-Pad2_ 0.75732k		

.end
