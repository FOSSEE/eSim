*noise of a resistive divider
*noise of a resistive divider with filter
*noise as above after a noiseless amplifier with gain 5

V1 1 0 dc 0 ac 1
R1 1 2 10k
R2 2 0 10k

V21 21 0 dc 0 ac 1
R21 21 22 10k
R22 22 0 10k
C22 22 0 1u

a1 2 3 amp
.model amp gain(in_offset = 0 gain = 5.0
+ out_offset = 0)

a2 22 23 amp

.control

noise v(2) V1 dec 10 1 100k
print onoise_total inoise_total
setplot noise1
print onoise_spectrum[0] inoise_spectrum[0]

noise v(3) V1 dec 10 1 100k
print onoise_total inoise_total
setplot noise3
print onoise_spectrum[0] inoise_spectrum[0]

noise v(22) V21 dec 10 1 100k
print onoise_total inoise_total
setplot noise5
print onoise_spectrum[0] inoise_spectrum[0]

noise v(23) V21 dec 10 1 100k
print onoise_total inoise_total
setplot noise7
print onoise_spectrum[0] inoise_spectrum[0]
set xbrushwidth = 2
plot  onoise_spectrum noise5.onoise_spectrum inoise_spectrum xlimit 1 1e5

.endc

.end


