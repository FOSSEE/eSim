* C:\Users\Bhargav\eSim\src\SubcircuitLibrary\4072\4072.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/31/19 10:17:30

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad5_ Net-_U1-Pad2_ Net-_U2-Pad3_ d_or		
U3  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U3-Pad3_ d_or		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ ? ? ? Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ ? PORT		
U4  Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U4-Pad3_ d_or		
U5  Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U5-Pad3_ d_or		
U6  Net-_U2-Pad3_ Net-_U3-Pad3_ Net-_U1-Pad1_ d_or		
U7  Net-_U4-Pad3_ Net-_U5-Pad3_ Net-_U1-Pad13_ d_or		

.end
