.title KiCad schematic
U1 unconnected-_U1-Pad1_ unconnected-_U1-Pad2_ unconnected-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ unconnected-_U1-Pad6_ unconnected-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT
U6 Net-_U1-Pad14_ Net-_U1-Pad14_ Net-_U2-Pad2_ unconnected-_U6-Pad4_ Net-_U5-Pad2_ Net-_U1-Pad9_ unconnected-_U6-Pad7_ d_jkff
U5 Net-_U11-Pad1_ Net-_U5-Pad2_ d_inverter
U2 Net-_U1-Pad10_ Net-_U2-Pad2_ d_inverter
U3 Net-_U1-Pad11_ Net-_U3-Pad2_ d_inverter
U7 Net-_U1-Pad14_ Net-_U1-Pad14_ Net-_U3-Pad2_ unconnected-_U7-Pad4_ Net-_U4-Pad2_ Net-_U1-Pad5_ unconnected-_U7-Pad7_ d_jkff
U4 Net-_U11-Pad1_ Net-_U4-Pad2_ d_inverter
U8 Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U11-Pad1_ d_nand
U13 Net-_U1-Pad14_ Net-_U1-Pad14_ Net-_U13-Pad3_ unconnected-_U13-Pad4_ Net-_U11-Pad2_ Net-_U1-Pad4_ unconnected-_U13-Pad7_ d_jkff
U9 Net-_U1-Pad5_ Net-_U13-Pad3_ d_inverter
U11 Net-_U11-Pad1_ Net-_U11-Pad2_ d_inverter
U12 Net-_U11-Pad1_ Net-_U12-Pad2_ d_inverter
U10 Net-_U1-Pad4_ Net-_U10-Pad2_ d_inverter
U14 Net-_U1-Pad14_ Net-_U1-Pad14_ Net-_U10-Pad2_ unconnected-_U14-Pad4_ Net-_U12-Pad2_ Net-_U1-Pad8_ unconnected-_U14-Pad7_ d_jkff
.end
