* C:\FOSSEE\eSim\library\SubcircuitLibrary\cmos_and\cmos_and.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/22/22 18:26:47

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_p		
M4  Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_p		
M2  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad4_ mosfet_n		
M3  Net-_M2-Pad3_ Net-_M3-Pad2_ Net-_M2-Pad4_ Net-_M2-Pad4_ mosfet_n		
U1  Net-_M1-Pad2_ Net-_M2-Pad4_ Net-_M1-Pad3_ Net-_M3-Pad2_ Net-_M5-Pad1_ PORT		
M6  Net-_M5-Pad1_ Net-_M1-Pad1_ Net-_M1-Pad3_ Net-_M1-Pad3_ mosfet_p		
M5  Net-_M5-Pad1_ Net-_M1-Pad1_ Net-_M2-Pad4_ Net-_M2-Pad4_ mosfet_n		

.end
