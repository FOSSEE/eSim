* /home/fossee/Downloads/eSim-master/Examples/CMOS_Inverter/CMOS_Inverter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Aug 19 14:20:52 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
C1  out 0 1u		
v1  in 0 dc		
v2  vcc 0 5		
M1  out in 0 0 MOS_N		
M2  out in vcc vcc MOS_P		

.end
