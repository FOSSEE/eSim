* C:\FOSSEE2\eSim\library\SubcircuitLibrary\LM113-PORT\LM113-PORT.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/18/24 10:50:46

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  Net-_R1-Pad1_ Net-_Q1-Pad2_ 200		
R2  Net-_R2-Pad1_ Net-_R1-Pad1_ 3.9k		
R3  Net-_R1-Pad1_ Net-_Q1-Pad1_ 170		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
R4  Net-_R2-Pad1_ Net-_C1-Pad2_ 13.5k		
Q2  Net-_C1-Pad2_ Net-_Q1-Pad1_ Net-_Q2-Pad3_ eSim_NPN		
R5  Net-_Q2-Pad3_ Net-_Q1-Pad3_ 1.6k		
R6  Net-_R2-Pad1_ Net-_Q4-Pad3_ 1.5k		
Q4  Net-_Q3-Pad1_ Net-_Q3-Pad1_ Net-_Q4-Pad3_ eSim_PNP		
Q3  Net-_Q3-Pad1_ Net-_Q1-Pad1_ Net-_Q3-Pad3_ eSim_NPN		
R7  Net-_Q3-Pad3_ Net-_Q1-Pad3_ 2k		
R8  Net-_R2-Pad1_ Net-_Q5-Pad3_ 1.5k		
Q5  Net-_C1-Pad1_ Net-_Q3-Pad1_ Net-_Q5-Pad3_ eSim_PNP		
Q6  Net-_C1-Pad1_ Net-_C1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
Q7  Net-_Q7-Pad1_ Net-_C1-Pad1_ Net-_C2-Pad1_ eSim_PNP		
R9  Net-_R2-Pad1_ Net-_C2-Pad1_ 10		
R10  Net-_C2-Pad2_ Net-_Q7-Pad1_ 3k		
Q8  Net-_Q7-Pad1_ Net-_Q1-Pad1_ Net-_Q8-Pad3_ eSim_NPN		
R11  Net-_Q8-Pad3_ Net-_Q1-Pad3_ 1.1k		
Q9  Net-_C2-Pad1_ Net-_Q7-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 75p		
C2  Net-_C2-Pad1_ Net-_C2-Pad2_ 30p		
U1  Net-_R2-Pad1_ Net-_Q1-Pad3_ PORT		

.end
