.title KiCad schematic
V_4B1 Net-_V_4B1-Pad1_ GND DC
U6 V_4Y plot_v1
U5 V_3Y plot_v1
U7 Net-_V_4B1-Pad1_ Net-_V_4A1-Pad1_ Net-_V_3B1-Pad1_ Net-_V_3A1-Pad1_ Net-_U7-Pad5_ Net-_U7-Pad6_ Net-_U7-Pad7_ Net-_U7-Pad8_ adc_bridge_4
v1 Net-_X1-Pad14_ GND 5
V_3A1 Net-_V_3A1-Pad1_ GND DC
V_3B1 Net-_V_3B1-Pad1_ GND DC
V_4A1 Net-_V_4A1-Pad1_ GND DC
U4 Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U4-Pad3_ Net-_U4-Pad4_ V_4Y V_3Y V_2Y V_1Y dac_bridge_4
U3 V_2Y plot_v1
V_2A1 Net-_V_2A1-Pad1_ GND DC
V_1B1 Net-_V_1B1-Pad1_ GND DC
V_1A1 Net-_V_1A1-Pad1_ GND DC
V_2B1 Net-_V_2B1-Pad1_ GND DC
X1 Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U4-Pad4_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U4-Pad3_ GND Net-_U4-Pad2_ Net-_U7-Pad8_ Net-_U7-Pad7_ Net-_U4-Pad1_ Net-_U7-Pad6_ Net-_U7-Pad5_ Net-_X1-Pad14_ 74HC86
U2 V_1Y plot_v1
U1 Net-_V_1A1-Pad1_ Net-_V_1B1-Pad1_ Net-_V_2A1-Pad1_ Net-_V_2B1-Pad1_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ adc_bridge_4
.end
