.title KiCad schematic
R9 GND Net-_Q10-Pad3_ 5k
R8 GND Net-_Q2-Pad1_ 2k
Q10 Net-_I4-Pad2_ Net-_I4-Pad2_ Net-_Q10-Pad3_ eSim_NPN
I5 Net-_I5-Pad1_ GND 500u
Q9 Net-_Q12-Pad2_ Net-_I4-Pad2_ Net-_Q2-Pad1_ eSim_NPN
Q4 Net-_Q4-Pad1_ vref Net-_I1-Pad1_ eSim_NPN
R3 vin Net-_I2-Pad1_ 1k
Q3 Net-_Q3-Pad1_ vref Net-_I2-Pad2_ eSim_PNP
Q2 Net-_Q2-Pad1_ vin Net-_I2-Pad2_ eSim_PNP
I2 Net-_I2-Pad1_ Net-_I2-Pad2_ 200u
R10 Net-_M1-Pad2_ Net-_I2-Pad1_ 10k
M1 Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_I2-Pad1_ Net-_I2-Pad1_ eSim_MOS_P
Q12 Net-_M4-Pad2_ Net-_Q12-Pad2_ Net-_I5-Pad1_ eSim_NPN
R11 Net-_M4-Pad2_ Net-_I2-Pad1_ 10k
Q11 Net-_M1-Pad2_ Net-_Q11-Pad2_ Net-_I5-Pad1_ eSim_NPN
M4 out Net-_M4-Pad2_ Net-_I2-Pad1_ Net-_I2-Pad1_ eSim_MOS_P
Q6 Net-_Q4-Pad1_ Net-_I3-Pad1_ Net-_Q11-Pad2_ eSim_PNP
R6 GND Net-_Q3-Pad1_ 2k
R5 Net-_Q4-Pad1_ Net-_I2-Pad1_ 50k
R4 Net-_Q5-Pad3_ Net-_I2-Pad1_ 50k
Q7 Net-_Q11-Pad2_ Net-_I4-Pad2_ Net-_Q3-Pad1_ eSim_NPN
Q5 Net-_I3-Pad1_ Net-_I3-Pad1_ Net-_Q5-Pad3_ eSim_PNP
I3 Net-_I3-Pad1_ GND 300u
M2 Net-_M1-Pad1_ Net-_M1-Pad1_ GND GND eSim_MOS_N
v1 Net-_I2-Pad1_ GND 5
M3 out Net-_M1-Pad1_ GND GND eSim_MOS_N
R7 Net-_Q1-Pad1_ Net-_I2-Pad1_ 20k
I4 Net-_I2-Pad1_ Net-_I4-Pad2_ 1m
Q8 Net-_Q1-Pad1_ Net-_I3-Pad1_ Net-_Q12-Pad2_ eSim_PNP
I1 Net-_I1-Pad1_ GND 400u
Q1 Net-_Q1-Pad1_ vin Net-_I1-Pad1_ eSim_NPN
R2 GND vref 1k
R1 vref Net-_I2-Pad1_ 3k
.end
