* C:\FOSSEE\eSim\library\SubcircuitLibrary\MC1489_0\MC1489_0.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/29/25 19:55:03

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  Net-_Q1-Pad1_ Net-_D1-Pad2_ Net-_D1-Pad1_ eSim_NPN		
Q2  Net-_Q2-Pad1_ Net-_Q1-Pad1_ Net-_D1-Pad1_ eSim_NPN		
Q3  Net-_Q3-Pad1_ Net-_Q2-Pad1_ Net-_D1-Pad1_ eSim_NPN		
R2  Net-_D1-Pad2_ Net-_D1-Pad1_ 10K		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
R5  Net-_R4-Pad1_ Net-_Q2-Pad1_ 5K		
R4  Net-_R4-Pad1_ Net-_Q1-Pad1_ 9K		
R6  Net-_R4-Pad1_ Net-_Q3-Pad1_ 1.7K		
R1  Net-_R1-Pad1_ Net-_D1-Pad2_ 3.8K		
R3  Net-_D1-Pad2_ Net-_Q1-Pad1_ 6.7K		
U1  Net-_R1-Pad1_ Net-_D1-Pad2_ Net-_R4-Pad1_ Net-_Q3-Pad1_ Net-_D1-Pad1_ PORT		

.end
