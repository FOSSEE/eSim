* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Jun 24 12:24:33 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
X1  8 7 6 2 half_adder		
X2  5 6 4 3 half_adder		
U1  8 7 5 4 1 PORT		
U2  3 2 1 d_or		

.end
