.title KiCad schematic
M4 Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M4-Pad3_ Net-_M1-Pad3_ eSim_MOS_N
v1 Net-_M1-Pad4_ GND 5
U1 Net-_U1-Pad1_ Net-_M1-Pad1_ Net-_M4-Pad3_ PORT
M5 Net-_M1-Pad1_ Net-_M5-Pad2_ Net-_M4-Pad3_ Net-_M1-Pad4_ eSim_MOS_P
M2 Net-_M1-Pad3_ Net-_M1-Pad2_ GND GND eSim_MOS_N
M3 Net-_M1-Pad1_ Net-_M3-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N
U6 Net-_U4-Pad2_ Net-_M3-Pad2_ dac_bridge_1
M1 Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad4_ eSim_MOS_P
U5 Net-_U2-Pad2_ Net-_M5-Pad2_ dac_bridge_1
U4 Net-_U2-Pad2_ Net-_U4-Pad2_ d_inverter
U3 Net-_U2-Pad2_ Net-_M1-Pad2_ dac_bridge_1
U2 Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter
.end
