* C:\Users\Shanthipriya\Desktop\madeeasy\FOSSEE\eSim\library\SubcircuitLibrary\74AC283\74AC283.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/07/25 22:10:48

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U6-Pad1_ Net-_X1-Pad5_ full_adder		
X2  Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_X1-Pad5_ Net-_U6-Pad2_ Net-_X2-Pad5_ full_adder		
X3  Net-_U4-Pad3_ Net-_U4-Pad4_ Net-_X2-Pad5_ Net-_U6-Pad3_ Net-_X3-Pad5_ full_adder		
X4  Net-_U5-Pad3_ Net-_U5-Pad4_ Net-_X3-Pad5_ Net-_U6-Pad4_ Net-_U6-Pad5_ full_adder		
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ adc_bridge_3		
U3  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U3-Pad3_ Net-_U3-Pad4_ adc_bridge_2		
U4  Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U4-Pad3_ Net-_U4-Pad4_ adc_bridge_2		
U5  Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U5-Pad3_ Net-_U5-Pad4_ adc_bridge_2		
U6  Net-_U6-Pad1_ Net-_U6-Pad2_ Net-_U6-Pad3_ Net-_U6-Pad4_ Net-_U6-Pad5_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ dac_bridge_5		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ ? ? PORT		

.end
