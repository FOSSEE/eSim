* H:\esim\eSim\library\SubcircuitLibrary\MUX_21\MUX_21.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/16/25 20:44:44

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__nfet_01v8		
SC2  Net-_SC1-Pad1_ Net-_SC2-Pad2_ Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__nfet_01v8		
U1  Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC2-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_SC1-Pad1_ PORT		
scmode1  SKY130mode		
X1  Net-_SC1-Pad2_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_SC2-Pad2_ CMOS_INVTR		

.end
