* C:\FOSSEE\eSim\library\SubcircuitLibrary\FCT827\FCT827.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/10/24 02:15:36

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U2-Pad2_ Net-_U3-Pad2_ Net-_U10-Pad2_ d_and		
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter		
U3  Net-_U1-Pad2_ Net-_U3-Pad2_ d_inverter		
U5  Net-_U1-Pad3_ Net-_U10-Pad2_ Net-_U1-Pad13_ d_tristate		
U6  Net-_U1-Pad4_ Net-_U10-Pad2_ Net-_U1-Pad14_ d_tristate		
U7  Net-_U1-Pad5_ Net-_U10-Pad2_ Net-_U1-Pad15_ d_tristate		
U8  Net-_U1-Pad6_ Net-_U10-Pad2_ Net-_U1-Pad16_ d_tristate		
U9  Net-_U1-Pad7_ Net-_U10-Pad2_ Net-_U1-Pad17_ d_tristate		
U10  Net-_U1-Pad8_ Net-_U10-Pad2_ Net-_U1-Pad18_ d_tristate		
U11  Net-_U1-Pad9_ Net-_U10-Pad2_ Net-_U1-Pad19_ d_tristate		
U12  Net-_U1-Pad10_ Net-_U10-Pad2_ Net-_U1-Pad20_ d_tristate		
U13  Net-_U1-Pad11_ Net-_U10-Pad2_ Net-_U1-Pad21_ d_tristate		
U14  Net-_U1-Pad12_ Net-_U10-Pad2_ Net-_U1-Pad22_ d_tristate		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U1-Pad18_ Net-_U1-Pad19_ Net-_U1-Pad20_ Net-_U1-Pad21_ Net-_U1-Pad22_ PORT		

.end
