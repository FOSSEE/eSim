* /home/saurabh/Desktop/eSim/Examples/Differentiator/Differentiator.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Fri Mar 27 17:56:03 2020

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  in GND pwl		
U1  in plot_v1		
U2  out plot_v1		
R1  in Net-_C1-Pad2_ 100k		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 10n		
R2  Net-_R2-Pad1_ GND 1k		
R3  Net-_C1-Pad1_ out 1k		
R4  out GND 1k		
X1  ? Net-_C1-Pad1_ Net-_R2-Pad1_ Net-_X1-Pad4_ ? out Net-_X1-Pad7_ ? lm_741		
v3  Net-_X1-Pad7_ GND DC		
v2  GND Net-_X1-Pad4_ DC		

.end
