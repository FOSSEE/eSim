* /home/fossee/eSim-Workspace/Diode_characteristics/Diode_characteristics.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Feb 23 16:11:16 2016

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  in GND DC		
D1  in out D		
R1  Net-_R1-Pad1_ GND 1k		
U1  out Net-_R1-Pad1_ plot_i2		

.end
