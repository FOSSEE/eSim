* /home/bhargav/eSim-Workspace/D_PULLUP_PULLDOWN_CHARACTERISTICS/D_PULLUP_PULLDOWN_CHARACTERISTICS.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jul  2 12:59:56 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  /1 d_pulldown		
U3  /1 Net-_U1-Pad1_ Net-_U3-Pad3_ d_and		
U4  Net-_U3-Pad3_ o dac_bridge_1		
U5  o plot_v1		
U1  Net-_U1-Pad1_ d_pullup		

.end
