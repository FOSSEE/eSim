* C:\Users\Aditya\eSim-Workspace\MC1455B_IC\MC1455B_IC.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/18/24 13:03:45

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R2  Out GND 1k		
R3  In Net-_R1-Pad1_ 5.1k		
C1  Net-_C1-Pad1_ GND 0.01u		
C2  Vcap GND 0.1u		
R1  Net-_R1-Pad1_ Vcap 100.9k		
v1  In GND DC		
X1  GND Vcap Out In Net-_C1-Pad1_ Vcap Net-_R1-Pad1_ In MC_1455B		
R4  In Out 1k		
U1  In plot_v1		
U2  Out plot_v1		
U3  Vcap plot_v1		

.end
