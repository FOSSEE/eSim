* C:\FOSSEE\eSim\library\SubcircuitLibrary\bidirectional_switch\bidirectional_switch.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/10/25 10:34:27

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M3-Pad3_ GND mosfet_n		
M4  Net-_M3-Pad1_ Net-_M4-Pad2_ Net-_M3-Pad3_ Net-_M4-Pad4_ mosfet_p		
U1  Net-_M3-Pad1_ Net-_M3-Pad3_ Net-_M3-Pad2_ PORT		
U3  Net-_M3-Pad2_ Net-_U2-Pad1_ adc_bridge_1		
U4  Net-_U2-Pad2_ Net-_M4-Pad2_ dac_bridge_1		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ d_inverter		
v1  Net-_M4-Pad4_ GND 5		

.end
