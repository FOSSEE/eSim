* C:\Users\senba\Desktop\FOSSEE\eSim\library\SubcircuitLibrary\74HC279\74HC279.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 12/17/25 11:27:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad1_ Net-_U2-Pad2_ d_inverter		
U3  Net-_U1-Pad2_ Net-_U3-Pad2_ d_inverter		
U4  Net-_U1-Pad3_ Net-_U4-Pad2_ d_inverter		
U5  Net-_U1-Pad4_ Net-_U10-Pad1_ d_inverter		
U6  Net-_U1-Pad5_ Net-_U11-Pad1_ d_inverter		
U7  Net-_U2-Pad2_ Net-_U14-Pad1_ d_inverter		
U8  Net-_U3-Pad2_ Net-_U8-Pad2_ d_inverter		
U9  Net-_U4-Pad2_ Net-_U9-Pad2_ d_inverter		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ d_inverter		
U11  Net-_U11-Pad1_ Net-_U11-Pad2_ d_inverter		
U14  Net-_U14-Pad1_ Net-_U14-Pad2_ Net-_U14-Pad3_ d_nand		
X1  Net-_U14-Pad3_ Net-_U8-Pad2_ Net-_U9-Pad2_ Net-_U14-Pad2_ 3_and		
U15  Net-_U14-Pad2_ Net-_U15-Pad2_ d_inverter		
U17  Net-_U15-Pad2_ Net-_U17-Pad2_ d_inverter		
U19  Net-_U17-Pad2_ Net-_U1-Pad6_ d_inverter		
U12  Net-_U10-Pad2_ Net-_U12-Pad2_ Net-_U12-Pad3_ d_nand		
U13  Net-_U12-Pad3_ Net-_U11-Pad2_ Net-_U12-Pad2_ d_nand		
U16  Net-_U12-Pad2_ Net-_U16-Pad2_ d_inverter		
U18  Net-_U16-Pad2_ Net-_U1-Pad7_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ PORT		

.end
