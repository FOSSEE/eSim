* C:\FOSSEE\eSim\library\SubcircuitLibrary\CD4015BC_edge\CD4015BC_edge.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 4/21/2025 9:52:10 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  da clka qa1 ra dff_edge		
X3  qa1 clka qa2 ra dff_edge		
X5  qa2 clka qa3 ra dff_edge		
X7  qa3 clka qa4 ra dff_edge		
X2  db clkb qb1 rb dff_edge		
X4  qb1 clkb qb2 rb dff_edge		
X6  qb2 clkb qb3 rb dff_edge		
X8  qb3 clkb qb4 rb dff_edge		

.end
