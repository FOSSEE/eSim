* C:\FOSSEE\eSim\library\SubcircuitLibrary\tl431_sub\tl431_sub.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 03/29/25 21:28:50

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad1_ /Anode eSim_NPN		
Q4  Net-_C1-Pad2_ Net-_Q2-Pad1_ Net-_Q4-Pad3_ eSim_NPN		
Q9  Net-_C2-Pad2_ Net-_Q9-Pad2_ /Anode eSim_NPN		
Q6  Net-_C1-Pad1_ Net-_C1-Pad2_ /Anode eSim_NPN		
R1  Net-_R1-Pad1_ Net-_Q2-Pad1_ 2.4k		
R3  Net-_R1-Pad1_ Net-_C1-Pad2_ 7.2k		
R4  Net-_Q4-Pad3_ /Anode 800		
R7  Net-_Q9-Pad2_ Net-_Q2-Pad1_ 1k		
R6  Net-_Q5-Pad3_ Net-_C1-Pad1_ 4k		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 20p		
Q5  Net-_Q5-Pad1_ Net-_Q1-Pad3_ Net-_Q5-Pad3_ eSim_NPN		
R2  Net-_Q1-Pad3_ Net-_R1-Pad1_ 3.28k		
Q1  /Cathode /Ref Net-_Q1-Pad3_ eSim_NPN		
Q3  Net-_C2-Pad2_ Net-_C2-Pad2_ /Ref eSim_NPN		
Q7  Net-_Q5-Pad1_ Net-_Q5-Pad1_ Net-_Q7-Pad3_ eSim_PNP		
Q8  Net-_C2-Pad2_ Net-_Q5-Pad1_ Net-_Q8-Pad3_ eSim_PNP		
R5  /Cathode Net-_Q7-Pad3_ 800		
R8  /Cathode Net-_Q8-Pad3_ 800		
D1  /Anode Net-_C2-Pad2_ eSim_Diode		
C2  /Cathode Net-_C2-Pad2_ 20p		
Q10  /Cathode Net-_C2-Pad2_ Net-_Q10-Pad3_ eSim_NPN		
R9  Net-_Q10-Pad3_ Net-_Q11-Pad2_ 150		
Q11  /Cathode Net-_Q11-Pad2_ /Anode eSim_NPN		
R10  /Anode Net-_Q11-Pad2_ 10k		
D2  /Anode /Cathode eSim_Diode		
U1  /Cathode /Ref /Anode PORT		

.end
