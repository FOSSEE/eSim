* C:\FOSSEE\eSim\library\SubcircuitLibrary\ic100117\ic100117.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/10/25 22:41:29

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U5  Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U5-Pad3_ d_or		
U6  Net-_U1-Pad24_ Net-_U1-Pad1_ Net-_U6-Pad3_ d_or		
X3  Net-_U5-Pad3_ Net-_U6-Pad3_ Net-_U1-Pad19_ Net-_U1-Pad4_ 3_and		
U9  Net-_U1-Pad4_ Net-_U1-Pad5_ d_inverter		
U10  Net-_U1-Pad22_ Net-_U1-Pad23_ Net-_U10-Pad3_ d_or		
U2  Net-_U1-Pad20_ Net-_U1-Pad21_ Net-_U2-Pad3_ d_or		
X1  Net-_U10-Pad3_ Net-_U2-Pad3_ Net-_U1-Pad17_ Net-_U1-Pad8_ 3_and		
U7  Net-_U1-Pad8_ Net-_U1-Pad9_ d_inverter		
U3  Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U3-Pad3_ d_or		
U4  Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U4-Pad3_ d_or		
X2  Net-_U3-Pad3_ Net-_U4-Pad3_ Net-_U1-Pad16_ Net-_U1-Pad11_ 3_and		
U8  Net-_U1-Pad11_ Net-_U1-Pad10_ d_inverter		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U1-Pad19_ Net-_U1-Pad20_ Net-_U1-Pad21_ Net-_U1-Pad22_ Net-_U1-Pad23_ Net-_U1-Pad24_ PORT		

.end
