* C:\FOSSEE\eSim\library\SubcircuitLibrary\mc1496\mc1496.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/12/25 22:39:35

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
Q5  Net-_Q5-Pad1_ Net-_Q5-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
Q6  Net-_Q2-Pad1_ Net-_Q5-Pad2_ Net-_Q6-Pad3_ eSim_NPN		
Q9  Net-_Q5-Pad1_ Net-_Q2-Pad2_ Net-_Q6-Pad3_ eSim_NPN		
Q3  Net-_Q2-Pad3_ Net-_Q3-Pad2_ Net-_Q3-Pad3_ eSim_NPN		
Q4  Net-_Q3-Pad3_ Net-_Q1-Pad1_ Net-_Q4-Pad3_ eSim_NPN		
Q7  Net-_Q6-Pad3_ Net-_Q7-Pad2_ Net-_Q7-Pad3_ eSim_NPN		
Q8  Net-_Q7-Pad3_ Net-_Q1-Pad1_ Net-_Q8-Pad3_ eSim_NPN		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad1_ Net-_Q1-Pad3_ eSim_NPN		
R2  Net-_Q4-Pad3_ Net-_R1-Pad2_ 500		
R1  Net-_Q1-Pad3_ Net-_R1-Pad2_ 500		
R3  Net-_Q8-Pad3_ Net-_R1-Pad2_ 500		
U1  Net-_Q7-Pad2_ Net-_Q7-Pad3_ Net-_Q3-Pad3_ Net-_Q3-Pad2_ Net-_Q1-Pad1_ Net-_Q2-Pad1_ ? Net-_Q2-Pad2_ ? Net-_Q5-Pad2_ ? Net-_Q5-Pad1_ ? Net-_R1-Pad2_ PORT		

.end
