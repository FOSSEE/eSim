* C:\Users\HP\OneDrive\Documents\FOSSEE\eSim\library\SubcircuitLibrary\TLC2201\TLC2201.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/15/25 15:12:39

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ /INV Net-_M1-Pad3_ /VDD mosfet_p		
M5  Net-_M1-Pad1_ /NON_INV Net-_C1-Pad1_ /VDD mosfet_p		
M2  Net-_M1-Pad3_ Net-_M1-Pad3_ /VSS /VSS mosfet_n		
M4  Net-_C1-Pad1_ Net-_M1-Pad3_ /VSS /VSS mosfet_n		
M3  /VDD Net-_M14-Pad2_ Net-_M1-Pad1_ /VDD mosfet_p		
M7  /VDD Net-_M14-Pad2_ Net-_M6-Pad1_ /VDD mosfet_p		
M10  /VDD Net-_M10-Pad2_ Net-_M10-Pad2_ /VDD mosfet_p		
M13  /VDD Net-_M10-Pad2_ /OUT /VDD mosfet_p		
M14  /VDD Net-_M14-Pad2_ Net-_M14-Pad2_ /VDD mosfet_p		
M17  /VDD Net-_M14-Pad2_ Net-_M15-Pad2_ /VDD mosfet_p		
M6  Net-_M6-Pad1_ Net-_C1-Pad1_ /VSS /VSS mosfet_n		
M8  Net-_M6-Pad1_ Net-_M6-Pad1_ /VSS /VSS mosfet_n		
M9  Net-_M10-Pad2_ Net-_M6-Pad1_ /VSS /VSS mosfet_n		
M12  /OUT Net-_C1-Pad1_ Net-_M11-Pad2_ /VSS mosfet_n		
M11  Net-_C1-Pad1_ Net-_M11-Pad2_ /VSS /VSS mosfet_n		
M15  Net-_M14-Pad2_ Net-_M15-Pad2_ Net-_M15-Pad3_ /VSS mosfet_n		
M16  Net-_M15-Pad2_ Net-_M15-Pad2_ Net-_D1-Pad1_ /VSS mosfet_n		
D1  Net-_D1-Pad1_ /VSS eSim_Diode		
R2  Net-_M15-Pad3_ /VSS 3k		
R1  Net-_M11-Pad2_ /VSS 3k		
C1  Net-_C1-Pad1_ /OUT 30p		
U1  ? /INV /NON_INV /VSS ? /VDD /OUT ? PORT		

.end
