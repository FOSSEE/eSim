* EESchema Netlist Version 1.1 (Spice format) creation date: Monday 17 December 2012 11:16:58 AM IST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  6 7 3 PORT		
Rout1  3 2 75		
Eout1  2 0 1 0 1		
Cbw1  1 0 31.85e-9		
Rbw1  1 4 0.5e6		
Ein1  4 0 7 6 100e3		
Rin1  7 6 2e6		

.end
