* eeschema netlist version 1.1 (spice format) creation date: 09/23/14 12:53:04
.include triac.sub
.include diac.sub

r3  1 2 250
c2  2 0 0.1u
* Plotting option vplot1
* Plotting option vplot1
x2  0 4 5 triac
x1  2 5 diac
c1  1 0 0.1u
r2  1 3 10k
v1  3 0 sine(0 100 50 0 0)
r1  4 3 100

.tran  10e-06 20e-03 0e-00
.plot v(2)
.plot v(3)
.plot v(3)-v(4) 
.end
