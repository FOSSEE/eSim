* /home/fossee/Downloads/eSim-master/Examples/rc/rc.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Aug 17 14:25:12 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  out in 1k		
C1  out GND 1u		
v1  in GND sine		

.end
