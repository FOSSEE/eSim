* E:\IC_74HC58\IC_74HC58.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/02/25 00:37:13

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U11-Pad6_ Net-_U11-Pad8_ Net-_U12-Pad7_ Net-_U12-Pad8_ Net-_U12-Pad9_ Net-_U12-Pad10_ Net-_U12-Pad11_ Net-_U12-Pad12_ Net-_U11-Pad5_ Net-_U11-Pad7_ Net-_U13-Pad1_ Net-_U14-Pad1_ 74HC58		
U12  A1 B1 C1 D1 E1 F1 Net-_U12-Pad7_ Net-_U12-Pad8_ Net-_U12-Pad9_ Net-_U12-Pad10_ Net-_U12-Pad11_ Net-_U12-Pad12_ adc_bridge_6		
U11  A2 B2 C2 D2 Net-_U11-Pad5_ Net-_U11-Pad6_ Net-_U11-Pad7_ Net-_U11-Pad8_ adc_bridge_4		
U13  Net-_U13-Pad1_ Y1 dac_bridge_1		
U14  Net-_U14-Pad1_ Y2 dac_bridge_1		
v1  A1 GND pulse		
v2  B1 GND pulse		
v3  C1 GND pulse		
v4  D1 GND pulse		
v5  E1 GND pulse		
v6  F1 GND pulse		
v7  A2 GND pulse		
v8  B2 GND pulse		
v9  C2 GND pulse		
v10  D2 GND pulse		
U15  Y1 plot_v1		
U16  Y2 plot_v1		
U1  A1 plot_v1		
U2  B1 plot_v1		
U3  C1 plot_v1		
U4  D1 plot_v1		
U5  E1 plot_v1		
U6  F1 plot_v1		
U7  A2 plot_v1		
U8  B2 plot_v1		
U9  C2 plot_v1		
U10  D2 plot_v1		

.end
