* D:\FOSSEE\eSim\library\SubcircuitLibrary\CA3045\CA3045.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/19/25 22:04:44

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_Q1-Pad3_ Net-_Q1-Pad2_ Net-_Q1-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ Net-_Q3-Pad2_ Net-_Q3-Pad1_ Net-_Q3-Pad3_ Net-_Q5-Pad2_ Net-_Q5-Pad1_ Net-_Q5-Pad3_ Net-_Q4-Pad2_ Net-_Q4-Pad1_ Net-_Q4-Pad3_ PORT		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ BC107		
Q2  Net-_Q1-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ BC107		
Q3  Net-_Q3-Pad1_ Net-_Q3-Pad2_ Net-_Q3-Pad3_ BC107		
Q5  Net-_Q5-Pad1_ Net-_Q5-Pad2_ Net-_Q5-Pad3_ BC107		
Q4  Net-_Q4-Pad1_ Net-_Q4-Pad2_ Net-_Q4-Pad3_ BC107		

.end
