* H:\esim\eSim\library\SubcircuitLibrary\Rnk_Blk\Rnk_Blk.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/17/25 16:26:27

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ PORT		
scmode1  SKY130mode		
X1  Net-_U1-Pad3_ Net-_U1-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_X1-Pad6_ DFF_CE		
X2  Net-_U1-Pad6_ Net-_X1-Pad6_ Net-_U1-Pad1_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_X2-Pad6_ MUX_21		
X3  Net-_U1-Pad3_ Net-_U1-Pad7_ Net-_X2-Pad6_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_X3-Pad6_ DFF_CE		
X4  Net-_U1-Pad8_ Net-_X3-Pad6_ Net-_X1-Pad6_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_X4-Pad6_ MUX_21		
X5  Net-_X4-Pad6_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad9_ Net-_U1-Pad10_ tri_state		

.end
