* C:\FOSSEE\eSim\library\SubcircuitLibrary\LT1460\LT1460.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/27/25 15:09:37

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R1  VOUT Net-_Q2-Pad2_ 150k		
R2  Net-_Q2-Pad2_ GND 48k		
Q2  Net-_Q1-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
Q4  Net-_Q3-Pad1_ Net-_Q2-Pad2_ Net-_Q4-Pad3_ eSim_NPN		
R5  Net-_Q4-Pad3_ Net-_Q2-Pad3_ 1k		
R6  Net-_Q2-Pad3_ GND 21k		
R3  VOUT Net-_Q1-Pad3_ 25k		
R4  VOUT Net-_Q3-Pad3_ 50k		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_PNP		
Q3  Net-_Q3-Pad1_ Net-_Q1-Pad2_ Net-_Q3-Pad3_ eSim_PNP		
Q5  GND Net-_Q3-Pad1_ Net-_Q1-Pad2_ eSim_PNP		
Q6  GND Net-_Q1-Pad1_ Net-_D1-Pad2_ eSim_PNP		
Q10  GND Net-_Q1-Pad1_ VOUT eSim_PNP		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q7  Net-_D1-Pad1_ Net-_Q7-Pad2_ VCC eSim_PNP		
Q8  Net-_Q7-Pad2_ Net-_Q7-Pad2_ VCC eSim_PNP		
Q9  Net-_Q7-Pad2_ Net-_D1-Pad1_ Net-_Q9-Pad3_ eSim_NPN		
R7  Net-_Q9-Pad3_ VOUT 100		
Q12  Net-_Q11-Pad1_ Net-_Q11-Pad1_ VCC eSim_PNP		
Q13  VOUT Net-_Q11-Pad1_ VCC eSim_PNP		
Q11  Net-_Q11-Pad1_ Net-_D1-Pad1_ VOUT eSim_NPN		
U1  VCC VOUT GND PORT		

.end
