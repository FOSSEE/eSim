* C:\FOSSEE\eSim\library\SubcircuitLibrary\bidirectional_shift_reg\bidirectional_shift_reg.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/02/25 13:59:38

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT		
U2  Net-_U2-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad8_ Net-_U1-Pad14_ dff_rst		
U5  Net-_U5-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad8_ Net-_U1-Pad13_ dff_rst		
U6  Net-_U6-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad8_ Net-_U1-Pad12_ dff_rst		
U8  Net-_U8-Pad1_ Net-_U1-Pad1_ Net-_U1-Pad8_ Net-_U1-Pad11_ dff_rst		
X4  Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U1-Pad12_ Net-_U1-Pad7_ Net-_U1-Pad2_ Net-_U1-Pad11_ Net-_U8-Pad1_ mux4		
X3  Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U1-Pad13_ Net-_U1-Pad11_ Net-_U1-Pad4_ Net-_U1-Pad12_ Net-_U6-Pad1_ mux4		
X2  Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U1-Pad14_ Net-_U1-Pad12_ Net-_U1-Pad5_ Net-_U1-Pad13_ Net-_U5-Pad1_ mux4		
X1  Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U1-Pad3_ Net-_U1-Pad13_ Net-_U1-Pad6_ Net-_U1-Pad14_ Net-_U2-Pad1_ mux4		

.end
