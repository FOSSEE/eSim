* /home/bhargav/eSim-Workspace/3_Input_NOR_Characteristics/3_Input_NOR_Characteristics.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Jul  2 12:47:46 2019

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U6  v1 v2 v3 Net-_U6-Pad4_ Net-_U6-Pad5_ Net-_U6-Pad6_ adc_bridge_3		
U10  v9 v8 v7 Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U10-Pad6_ adc_bridge_3		
v3  v1 GND DC		
v4  v2 GND DC		
v5  v3 GND DC		
U3  v1 plot_v1		
U4  v2 plot_v1		
U5  v3 plot_v1		
v1  v4 GND DC		
v2  v5 GND DC		
U1  v4 plot_v1		
U2  v5 plot_v1		
v6  v6 GND DC		
U14  v6 plot_v1		
v7  v7 GND DC		
v8  v8 GND DC		
v9  v9 GND DC		
U15  v7 plot_v1		
U16  v8 plot_v1		
U17  v9 plot_v1		
U8  Net-_U8-Pad1_ Net-_U8-Pad2_ Net-_U8-Pad3_ o1 o2 o3 dac_bridge_3		
U7  v4 v5 Net-_U7-Pad3_ Net-_U7-Pad4_ adc_bridge_2		
U11  v6 Net-_U11-Pad2_ adc_bridge_1		
U9  o1 plot_v1		
U12  o2 plot_v1		
U13  o3 plot_v1		
X1  Net-_U7-Pad3_ Net-_U7-Pad4_ Net-_U6-Pad4_ Net-_U6-Pad5_ Net-_U6-Pad6_ Net-_U8-Pad1_ ? Net-_U11-Pad2_ Net-_U8-Pad2_ Net-_U8-Pad3_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U10-Pad6_ ? IC_4025		

.end
