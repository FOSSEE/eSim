.title KiCad schematic
Q11 Net-_Q11-Pad1_ Net-_Q10-Pad1_ GND eSim_NPN
U1 Net-_D1-Pad1_ Net-_D4-Pad1_ Net-_Q11-Pad1_ PORT
Q7 Net-_Q7-Pad1_ Net-_Q10-Pad2_ GND eSim_NPN
Q9 Net-_Q10-Pad1_ Net-_Q11-Pad1_ Net-_Q7-Pad1_ eSim_PNP
Q10 Net-_Q10-Pad1_ Net-_Q10-Pad2_ GND eSim_NPN
Q8 Net-_Q11-Pad1_ Net-_Q7-Pad1_ Net-_Q10-Pad1_ eSim_NPN
I3 Net-_I1-Pad1_ Net-_D3-Pad1_ 0.2u
I4 Net-_I1-Pad1_ Net-_Q7-Pad1_ 6u
D2 Net-_D2-Pad1_ Net-_D1-Pad2_ eSim_Diode
I1 Net-_I1-Pad1_ Net-_D2-Pad1_ 0.2u
I2 Net-_I1-Pad1_ Net-_Q2-Pad3_ 5u
Q2 Net-_Q2-Pad1_ Net-_D1-Pad2_ Net-_Q2-Pad3_ eSim_PNP
Q1 GND Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_PNP
D1 Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode
D3 Net-_D3-Pad1_ Net-_D3-Pad2_ eSim_Diode
D4 Net-_D4-Pad1_ Net-_D3-Pad2_ eSim_Diode
Q6 GND Net-_D4-Pad1_ Net-_D3-Pad2_ eSim_PNP
Q4 Net-_Q10-Pad2_ Net-_Q2-Pad1_ GND eSim_NPN
Q5 Net-_Q10-Pad2_ Net-_D3-Pad2_ Net-_Q2-Pad3_ eSim_PNP
Q3 Net-_Q2-Pad1_ Net-_Q2-Pad1_ GND eSim_NPN
.end
