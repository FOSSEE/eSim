* C:\FOSSEE\eSim\library\SubcircuitLibrary\LT1004\LT1004.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 04/24/25 16:48:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q1  cathode Net-_C1-Pad1_ anode eSim_NPN		
Q2  Net-_C1-Pad1_ Net-_C1-Pad2_ cathode eSim_PNP		
R1  Net-_C1-Pad1_ anode 500k		
R2  cathode Net-_Q3-Pad3_ 7.5k		
Q3  Net-_C1-Pad2_ Net-_C1-Pad2_ Net-_Q3-Pad3_ eSim_PNP		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 20p		
Q4  Net-_C1-Pad2_ Net-_C2-Pad1_ Net-_Q4-Pad3_ eSim_NPN		
R3  Net-_Q4-Pad3_ anode 500		
Q5  Net-_C2-Pad1_ Net-_C2-Pad2_ cathode eSim_PNP		
Q6  Net-_C2-Pad1_ Net-_Q10-Pad2_ Net-_Q6-Pad3_ eSim_NPN		
R4  Net-_Q6-Pad3_ anode 60k		
R5  cathode Net-_Q10-Pad2_ 600k		
Q7  Net-_Q10-Pad2_ Net-_Q10-Pad2_ anode eSim_NPN		
Q8  Net-_C2-Pad2_ Net-_Q11-Pad1_ cathode eSim_PNP		
Q9  Net-_C2-Pad2_ Net-_Q9-Pad2_ Net-_Q10-Pad1_ eSim_NPN		
C2  Net-_C2-Pad1_ Net-_C2-Pad2_ 20p		
Q11  Net-_Q11-Pad1_ Net-_Q11-Pad1_ cathode eSim_PNP		
Q12  Net-_Q11-Pad1_ Net-_Q12-Pad2_ Net-_Q10-Pad1_ eSim_NPN		
Q10  Net-_Q10-Pad1_ Net-_Q10-Pad2_ anode eSim_NPN		
R6  cathode Net-_Q9-Pad2_ 200k		
R7  Net-_Q9-Pad2_ Net-_Q12-Pad2_ 50k		
R8  Net-_Q12-Pad2_ Net-_Q13-Pad3_ 300k		
Q13  anode anode Net-_Q13-Pad3_ eSim_PNP		
U1  cathode anode PORT		

.end
