* C:\FOSSEE\eSim\library\SubcircuitLibrary\74LVC1G17\74LVC1G17.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/16/26 00:21:49

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M4  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M3-Pad1_ VDD eSim_MOS_P		
M3  Net-_M3-Pad1_ Net-_M1-Pad2_ VDD VDD eSim_MOS_P		
M5  GND Net-_M1-Pad1_ Net-_M3-Pad1_ VDD eSim_MOS_P		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ GND eSim_MOS_N		
M2  Net-_M1-Pad3_ Net-_M1-Pad2_ GND GND eSim_MOS_N		
M6  VDD Net-_M1-Pad1_ Net-_M1-Pad3_ GND eSim_MOS_N		
M10  Net-_M10-Pad1_ Net-_M1-Pad1_ Net-_M10-Pad3_ VDD eSim_MOS_P		
M9  Net-_M10-Pad3_ Net-_M1-Pad1_ VDD VDD eSim_MOS_P		
M11  GND Net-_M10-Pad1_ Net-_M10-Pad3_ VDD eSim_MOS_P		
M7  Net-_M10-Pad1_ Net-_M1-Pad1_ Net-_M12-Pad3_ GND eSim_MOS_N		
M8  Net-_M12-Pad3_ Net-_M1-Pad1_ GND GND eSim_MOS_N		
M12  VDD Net-_M10-Pad1_ Net-_M12-Pad3_ GND eSim_MOS_N		
U1  Net-_M1-Pad2_ GND VDD Net-_M10-Pad1_ PORT		

.end
