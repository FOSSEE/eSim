.title KiCad schematic
Q3 Net-_Q1-Pad2_ Net-_Q3-Pad2_ Net-_Q1-Pad3_ eSim_NPN
Q1 Net-_C1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN
Q6 Net-_Q3-Pad2_ Net-_Q3-Pad2_ Net-_Q1-Pad3_ eSim_NPN
Q5 Net-_C2-Pad2_ Net-_Q5-Pad2_ Net-_Q3-Pad2_ eSim_NPN
Q8 Net-_Q5-Pad2_ Net-_Q5-Pad2_ Net-_Q3-Pad2_ eSim_NPN
Q10 Net-_Q10-Pad1_ Net-_Q10-Pad2_ Net-_Q1-Pad3_ eSim_NPN
Q9 Net-_Q12-Pad2_ Net-_Q12-Pad2_ Net-_Q10-Pad1_ eSim_NPN
Q12 Net-_Q11-Pad2_ Net-_Q12-Pad2_ Net-_Q10-Pad2_ eSim_NPN
R7 Net-_Q17-Pad2_ Net-_C1-Pad1_ 15.6k
U1 Net-_C1-Pad1_ Net-_R10-Pad2_ Net-_Q1-Pad3_ PORT
R6 Net-_C2-Pad1_ Net-_C1-Pad1_ 49k
R4 Net-_Q16-Pad1_ Net-_C1-Pad1_ 49k
Q17 Net-_C2-Pad1_ Net-_Q17-Pad2_ Net-_Q15-Pad1_ eSim_NPN
Q16 Net-_Q16-Pad1_ Net-_Q16-Pad2_ Net-_Q15-Pad1_ eSim_NPN
Q14 Net-_Q11-Pad2_ Net-_Q11-Pad2_ Net-_C1-Pad1_ eSim_PNP
R8 Net-_Q16-Pad2_ Net-_Q17-Pad2_ 600
R5 Net-_Q1-Pad3_ Net-_Q15-Pad3_ 1.1k
Q15 Net-_Q15-Pad1_ Net-_Q10-Pad1_ Net-_Q15-Pad3_ eSim_NPN
R9 Net-_Q1-Pad3_ Net-_Q16-Pad2_ 13.8k
R10 Net-_Q16-Pad2_ Net-_R10-Pad2_ 10k
Q13 Net-_Q10-Pad2_ Net-_Q10-Pad1_ Net-_Q13-Pad3_ eSim_NPN
R3 Net-_Q1-Pad3_ Net-_Q13-Pad3_ 2k
Q2 Net-_C1-Pad1_ Net-_C2-Pad2_ Net-_Q1-Pad2_ eSim_NPN
C1 Net-_C1-Pad1_ Net-_C1-Pad2_ 3pf
R1 Net-_C1-Pad2_ Net-_C2-Pad2_ 10k
Q4 Net-_C2-Pad2_ Net-_C2-Pad1_ Net-_Q11-Pad1_ eSim_PNP
R2 Net-_Q12-Pad2_ Net-_C1-Pad1_ 50k
Q11 Net-_Q11-Pad1_ Net-_Q11-Pad2_ Net-_C1-Pad1_ eSim_PNP
C2 Net-_C2-Pad1_ Net-_C2-Pad2_ 3pf
Q7 Net-_Q5-Pad2_ Net-_Q16-Pad1_ Net-_Q11-Pad1_ eSim_PNP
.end
