* H:\esim\eSim\library\SubcircuitLibrary\CMOS_INVTR\CMOS_INVTR.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 07/12/25 16:02:08

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad3_ sky130_fd_pr__pfet_01v8		
SC2  Net-_SC1-Pad1_ Net-_SC1-Pad2_ Net-_SC2-Pad3_ Net-_SC2-Pad3_ sky130_fd_pr__nfet_01v8		
U1  Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC2-Pad3_ Net-_SC1-Pad1_ PORT		
scmode1  SKY130mode		

.end
