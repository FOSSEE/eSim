* C:\Users\pavithra\eSim-Workspace\MC14076B_test\MC14076B_test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/20/25 17:49:07

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U6  Net-_U6-Pad1_ Net-_U6-Pad2_ Net-_U6-Pad3_ Net-_U6-Pad4_ adc_bridge_2		
v1  Net-_U6-Pad1_ GND DC		
v3  Net-_U6-Pad2_ GND DC		
U8  Net-_U8-Pad1_ Net-_U8-Pad2_ Net-_U8-Pad3_ Net-_U8-Pad4_ W X Y Z dac_bridge_4		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U10-Pad4_ adc_bridge_2		
v6  Net-_U10-Pad1_ GND DC		
v5  Net-_U10-Pad2_ GND DC		
U11  RST A B C D Net-_U11-Pad6_ Net-_U11-Pad7_ Net-_U11-Pad8_ Net-_U11-Pad9_ Net-_U11-Pad10_ adc_bridge_5		
v7  D GND pulse		
v8  C GND pulse		
v9  B GND pulse		
v10  A GND pulse		
v11  RST GND pulse		
U9  Net-_U9-Pad1_ Net-_U9-Pad2_ adc_bridge_1		
v4  Net-_U9-Pad1_ GND DC		
U4  W plot_v1		
U2  X plot_v1		
U1  Y plot_v1		
U3  Z plot_v1		
U7  CLK Net-_U7-Pad2_ adc_bridge_1		
v2  CLK GND pulse		
U5  CLK plot_v1		
U12  RST plot_v1		
U13  A plot_v1		
U14  B plot_v1		
U15  C plot_v1		
U16  D plot_v1		
X1  Net-_U6-Pad3_ Net-_U6-Pad4_ Net-_U8-Pad1_ Net-_U8-Pad2_ Net-_U8-Pad3_ Net-_U8-Pad4_ Net-_U7-Pad2_ GND Net-_U10-Pad4_ Net-_U10-Pad3_ Net-_U11-Pad10_ Net-_U11-Pad9_ Net-_U11-Pad8_ Net-_U11-Pad7_ Net-_U11-Pad6_ Net-_U9-Pad2_ MC14076B		

.end
