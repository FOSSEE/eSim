* C:\FOSSEE\eSim\library\SubcircuitLibrary\74V1G14\74V1G14.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 8/3/2022 1:17:12 AM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  /Vout /Inp Net-_M1-Pad3_ /GND mosfet_n		
M2  Net-_M1-Pad3_ /Inp /GND /GND mosfet_n		
M3  /Vcc /Inp Net-_M3-Pad3_ /Vcc mosfet_p		
M4  Net-_M3-Pad3_ /Inp /Vout /Vcc mosfet_p		
M5  /GND /Vout Net-_M3-Pad3_ /Vcc mosfet_p		
M6  /Vcc /Vout Net-_M1-Pad3_ /GND mosfet_n		
U1  ? /Inp /GND /Vout /Vcc PORT		

.end
