* C:\FOSSEE\eSim\library\SubcircuitLibrary\mc1489A\mc1489A.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/09/25 01:17:36

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ gnd Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ PORT		
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad14_ Net-_U1-Pad3_ gnd MC1489A_0		
X3  Net-_U1-Pad10_ Net-_U1-Pad9_ Net-_U1-Pad14_ Net-_U1-Pad8_ gnd MC1489A_0		
X2  Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad14_ Net-_U1-Pad6_ gnd MC1489A_0		
X4  Net-_U1-Pad13_ Net-_U1-Pad12_ Net-_U1-Pad14_ Net-_U1-Pad11_ gnd MC1489A_0		

.end
