.title KiCad schematic
U4 Net-_U2-Pad3_ Net-_U3-Pad3_ Net-_U4-Pad3_ d_and
U1 Net-_U1-Pad1_ Net-_U1-Pad2_ unconnected-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ unconnected-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ unconnected-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ unconnected-_U1-Pad14_ PORT
U2 Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad3_ d_and
U3 Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U3-Pad3_ d_and
U5 Net-_U4-Pad3_ Net-_U1-Pad6_ d_inverter
U9 Net-_U8-Pad3_ Net-_U1-Pad8_ d_inverter
U8 Net-_U6-Pad3_ Net-_U7-Pad3_ Net-_U8-Pad3_ d_and
U6 Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U6-Pad3_ d_and
U7 Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U7-Pad3_ d_and
.end
