* C:\Users\Aditya\eSim-Workspace\CA3240_IC_Test\CA3240_IC_Test.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/26/24 18:38:14

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_C1-Pad1_ Net-_C1-Pad2_ Net-_R3-Pad2_ Net-_X1-Pad4_ Net-_X1-Pad5_ Net-_C2-Pad2_ Net-_C2-Pad1_ Net-_R5-Pad1_ C3240_IC		
v3  Net-_X1-Pad5_ GND DC		
v1  Vin1 GND sine		
R3  Vin1 Net-_R3-Pad2_ 1000k		
R2  Net-_C1-Pad2_ Net-_C1-Pad1_ 100k		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 2000p		
R1  Net-_R1-Pad1_ Net-_C1-Pad2_ 10k		
R4  Net-_R1-Pad1_ Net-_C2-Pad1_ 10k		
R6  Net-_C2-Pad2_ Net-_C2-Pad1_ 100k		
C2  Net-_C2-Pad1_ Net-_C2-Pad2_ 2000p		
R5  Net-_R5-Pad1_ Vin2 1000k		
v4  Vin2 GND sine		
v2  Net-_X1-Pad4_ GND DC		
X2  Vout Net-_R10-Pad2_ Net-_R11-Pad2_ Net-_X2-Pad4_ Net-_X2-Pad5_ ? ? ? C3240_IC		
v5  Net-_X2-Pad4_ GND DC		
v6  Net-_X2-Pad5_ GND DC		
R8  Net-_R11-Pad2_ Net-_C1-Pad1_ 100k		
R7  Net-_R10-Pad2_ Net-_C2-Pad2_ 100k		
R9  Vout GND 10k		
U1  Vin1 plot_v1		
U2  Vin2 plot_v1		
U3  Vout plot_v1		
R10  Vout Net-_R10-Pad2_ 100k		
R11  GND Net-_R11-Pad2_ 100k		

.end
