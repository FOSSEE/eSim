* C:\FOSSEE\eSim\library\SubcircuitLibrary\Buffer\Buffer.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/28/24 23:00:30

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_U1-Pad1_ Net-_X1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ NOT_Gate		
X2  Net-_X1-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ NOT_Gate		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ PORT		

.end
