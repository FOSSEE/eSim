* EESchema Netlist Version 1.1 (Spice format) creation date: Thu May  7 15:36:48 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U3  4 5 19 12 28 9 25 d_jkff		
v1  2 20 dc		
v3  1 20 dc		
v4  33 20 0		
v2  3 20 pulse		
U5  25 25 19 11 29 21 34 d_jkff		
U7  35 35 19 17 30 22 36 d_jkff		
U10  27 27 19 18 16 23 20 d_jkff		
U6  34 25 35 d_and		
U8  36 35 27 d_and		
U4  26 33 31 32 28 29 30 16 adc_bridge_4		
v10  31 20 0		
v11  32 20 0		
v9  26 20 0		
v8  14 20 0		
U2  15 14 10 13 18 17 11 12 adc_bridge_4		
v6  10 20 0		
v7  13 20 0		
v5  15 20 0		
U1  2 3 1 4 19 5 adc_bridge_3		
U9  9 21 22 23 6 7 8 24 dac_bridge_4		
R2  20 7 1k		
R3  20 8 1k		
R4  20 24 1k		
R1  20 6 1k		

.end
