* C:\Users\HP\OneDrive\Documents\FOSSEE\eSim\library\SubcircuitLibrary\8286\8286.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 05/22/25 01:06:17

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  /OE_BAR /TRANS/RXR_BAR Net-_U11-Pad2_ d_nor		
U2  /TRANS/RXR_BAR Net-_U2-Pad2_ d_inverter		
U6  /A0 Net-_U10-Pad2_ /B0 d_tristate		
U8  /A1 Net-_U10-Pad2_ /B1 d_tristate		
U10  /A2 Net-_U10-Pad2_ /B2 d_tristate		
U16  /A4 Net-_U10-Pad2_ /B4 d_tristate		
U18  /A5 Net-_U10-Pad2_ /B5 d_tristate		
U20  /A6 Net-_U10-Pad2_ /B6 d_tristate		
U22  /A7 Net-_U10-Pad2_ /B7 d_tristate		
U5  /B0 Net-_U11-Pad2_ /A0 d_tristate		
U7  /B1 Net-_U11-Pad2_ /A1 d_tristate		
U9  /B2 Net-_U11-Pad2_ /A2 d_tristate		
U15  /B4 Net-_U11-Pad2_ /A4 d_tristate		
U17  /B5 Net-_U11-Pad2_ /A5 d_tristate		
U19  /B6 Net-_U11-Pad2_ /A6 d_tristate		
U21  /B7 Net-_U11-Pad2_ /A7 d_tristate		
U1  /OE_BAR /TRANS/RXR_BAR /A0 /B0 /A1 /B1 /A2 /B2 /A3 /B3 /A4 /B4 /A5 /B5 /A6 /B6 /A7 /B7 ? ? PORT		
U11  /B3 Net-_U11-Pad2_ /A3 d_tristate		
U12  /A3 Net-_U10-Pad2_ /B3 d_tristate		
U4  Net-_U2-Pad2_ /OE_BAR Net-_U10-Pad2_ d_nor		

.end
