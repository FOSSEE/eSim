* C:\FOSSEE\eSim\library\SubcircuitLibrary\AND_3\AND_3.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/05/24 11:17:24

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M3  Net-_M1-Pad3_ Net-_M1-Pad2_ Net-_M3-Pad3_ Net-_M3-Pad3_ mosfet_n		
M4  Net-_M3-Pad3_ Net-_M2-Pad2_ Net-_M4-Pad3_ Net-_M4-Pad3_ mosfet_n		
M5  Net-_M4-Pad3_ Net-_M5-Pad2_ Net-_M5-Pad3_ Net-_M5-Pad3_ mosfet_n		
M7  Net-_M7-Pad1_ Net-_M1-Pad3_ Net-_M5-Pad3_ Net-_M5-Pad3_ mosfet_n		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M2  Net-_M1-Pad1_ Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M6  Net-_M1-Pad1_ Net-_M5-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad1_ mosfet_p		
M8  Net-_M1-Pad1_ Net-_M1-Pad3_ Net-_M7-Pad1_ Net-_M1-Pad1_ mosfet_p		
U1  Net-_M1-Pad2_ Net-_M2-Pad2_ Net-_M5-Pad2_ Net-_M5-Pad3_ Net-_M1-Pad1_ Net-_M7-Pad1_ PORT		

.end
