* C:\FOSSEE\eSim\library\SubcircuitLibrary\AD744_Subcircuit\AD744_Subcircuit.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 02/02/25 20:54:37

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
I1  Net-_I1-Pad1_ Net-_I1-Pad2_ 400uA		
R1  Net-_I1-Pad1_ Net-_Q1-Pad1_ 300		
R3  Net-_I1-Pad1_ Net-_Q3-Pad1_ 300		
R2  Net-_D1-Pad2_ Net-_Q5-Pad3_ 1k		
Q2  Net-_Q2-Pad1_ Net-_Q2-Pad2_ Net-_Q2-Pad3_ eSim_NPN		
R4  Net-_Q2-Pad3_ Net-_Q5-Pad3_ 1k		
Q4  Net-_I1-Pad2_ Net-_Q2-Pad1_ Net-_Q4-Pad3_ eSim_NPN		
C1  Net-_C1-Pad1_ Net-_C1-Pad2_ 5pF		
Q5  Net-_C1-Pad1_ Net-_Q4-Pad3_ Net-_Q5-Pad3_ eSim_NPN		
R5  Net-_Q4-Pad3_ Net-_Q5-Pad3_ 8k		
I2  Net-_D2-Pad1_ Net-_I1-Pad2_ 2mA		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
D2  Net-_D2-Pad1_ Net-_D2-Pad2_ eSim_Diode		
D3  Net-_D2-Pad2_ Net-_C1-Pad1_ eSim_Diode		
Q7  Net-_Q5-Pad3_ Net-_C1-Pad1_ Net-_Q6-Pad3_ eSim_PNP		
Q6  Net-_I1-Pad2_ Net-_D2-Pad1_ Net-_Q6-Pad3_ eSim_NPN		
U1  Net-_Q1-Pad2_ Net-_C1-Pad2_ Net-_Q2-Pad2_ Net-_Q3-Pad2_ Net-_I1-Pad2_ Net-_Q6-Pad3_ Net-_C1-Pad1_ Net-_Q5-Pad3_ PORT		
Q3  Net-_Q3-Pad1_ Net-_Q3-Pad2_ Net-_Q2-Pad1_ eSim_NPN		
Q1  Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_D1-Pad1_ eSim_NPN		

.end
