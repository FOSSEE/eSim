* C:\FOSSEE\eSim\library\SubcircuitLibrary\cd4070b_ic\cd4070b_ic.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/23/25 22:05:51

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M3  Net-_M11-Pad1_ Net-_M1-Pad2_ Net-_M1-Pad1_ Net-_M11-Pad1_ eSim_MOS_P		
M2  Net-_M2-Pad1_ Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
M4  Net-_M11-Pad1_ Net-_M2-Pad2_ Net-_M2-Pad1_ Net-_M11-Pad1_ eSim_MOS_P		
M6  Net-_M1-Pad1_ Net-_M2-Pad2_ Net-_M10-Pad2_ Net-_M11-Pad1_ eSim_MOS_P		
M5  Net-_M1-Pad1_ Net-_M2-Pad1_ Net-_M10-Pad2_ Net-_M1-Pad3_ eSim_MOS_N		
M8  Net-_M11-Pad1_ Net-_M2-Pad1_ Net-_M8-Pad3_ Net-_M11-Pad1_ eSim_MOS_P		
M9  Net-_M8-Pad3_ Net-_M1-Pad1_ Net-_M10-Pad2_ Net-_M11-Pad1_ eSim_MOS_P		
M7  Net-_M10-Pad2_ Net-_M1-Pad1_ Net-_M2-Pad1_ Net-_M1-Pad3_ eSim_MOS_N		
M11  Net-_M11-Pad1_ Net-_M10-Pad2_ Net-_M10-Pad1_ Net-_M11-Pad1_ eSim_MOS_P		
M10  Net-_M10-Pad1_ Net-_M10-Pad2_ Net-_M1-Pad3_ Net-_M1-Pad3_ eSim_MOS_N		
U1  Net-_M2-Pad2_ Net-_M1-Pad2_ Net-_M10-Pad1_ Net-_M10-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad2_ Net-_M1-Pad3_ Net-_M2-Pad2_ Net-_M1-Pad2_ Net-_M10-Pad1_ Net-_M10-Pad1_ Net-_M1-Pad2_ Net-_M2-Pad2_ Net-_M11-Pad1_ PORT		

.end
