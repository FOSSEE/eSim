* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/SN54L98/SN54L98.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Jul 10 12:28:04 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X2  Net-_U1-Pad5_ Net-_X1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad6_ Net-_U1-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad13_ DS_blk		
X3  Net-_U1-Pad7_ Net-_X1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad8_ Net-_U1-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad14_ DS_blk		
X4  Net-_U1-Pad9_ Net-_X1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad10_ Net-_U1-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad15_ DS_blk		
X5  Net-_U1-Pad11_ Net-_X1-Pad4_ Net-_U1-Pad1_ Net-_U1-Pad12_ Net-_U1-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad16_ DS_blk		
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_X1-Pad4_ CMOS_INVTR		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ PORT		
scmode1  SKY130mode		

.end
