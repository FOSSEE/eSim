* /home/fossee/Downloads/eSim-master/Examples/Inverting_Amplifier/Inverting_Amplifier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Wed Aug 19 15:19:14 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_R2-Pad2_ Net-_R1-Pad2_ Out UA741		
v1  In GND sine		
R2  GND Net-_R2-Pad2_ 1k		
R1  In Net-_R1-Pad2_ 1k		
R5  Net-_R1-Pad2_ Out 2k		
R3  Out GND 1k		

.end
