* C:\Users\Aditya\eSim-Workspace\SN74F521\SN74F521.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 08/24/24 18:28:18

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
x1  OE_BAR P0 Q0 P1 Q1 P2 Q2 P3 Q3 GND P4 Q4 P5 Q5 P6 Q6 P7 Q7 OUT Net-_v2-Pad1_ SN74F521_IC		
v1  P0 GND pulse		
v2  Net-_v2-Pad1_ GND DC		
R2  OUT GND 1000k		
R1  GND OE_BAR 1000k		
U2  OUT plot_v1		
U1  OE_BAR plot_v1		
v3  Q0 GND pulse		
v4  P1 GND pulse		
v5  Q1 GND pulse		
v6  P2 GND pulse		
v7  Q2 GND pulse		
v8  P3 GND pulse		
v9  Q3 GND pulse		
v10  P4 GND pulse		
v11  Q4 GND pulse		
v12  P5 GND pulse		
v13  Q5 GND pulse		
v14  P6 GND pulse		
v15  Q6 GND pulse		
v16  P7 GND pulse		
v17  Q7 GND pulse		
U18  Q7 plot_v1		
U17  P7 plot_v1		
U16  Q6 plot_v1		
U15  P6 plot_v1		
U14  Q5 plot_v1		
U13  P5 plot_v1		
U12  Q4 plot_v1		
U11  P4 plot_v1		
U10  Q3 plot_v1		
U9  P3 plot_v1		
U8  Q2 plot_v1		
U7  P2 plot_v1		
U6  Q1 plot_v1		
U5  P1 plot_v1		
U4  Q0 plot_v1		
U3  P0 plot_v1		

.end
