.title KiCad schematic
U1 Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ GND Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ GND PORT
U6 Net-_U1-Pad15_ Net-_X5-Pad4_ d_inverter
X2 Net-_X1-Pad1_ Net-_U2-Pad2_ Net-_U5-Pad2_ Net-_U1-Pad5_ Net-_X2-Pad5_ 4_and
X1 Net-_X1-Pad1_ Net-_U2-Pad2_ Net-_U3-Pad2_ Net-_U1-Pad6_ Net-_X1-Pad5_ 4_and
X3 Net-_X1-Pad1_ Net-_U4-Pad2_ Net-_U3-Pad2_ Net-_U1-Pad4_ Net-_X3-Pad5_ 4_and
U4 Net-_U2-Pad2_ Net-_U4-Pad2_ d_inverter
U5 Net-_U3-Pad2_ Net-_U5-Pad2_ d_inverter
U2 Net-_U1-Pad2_ Net-_U2-Pad2_ d_inverter
U3 Net-_U1-Pad14_ Net-_U3-Pad2_ d_inverter
X9 Net-_X1-Pad5_ Net-_X2-Pad5_ Net-_X3-Pad5_ Net-_X4-Pad5_ Net-_U1-Pad7_ 4_OR
X6 Net-_U1-Pad11_ Net-_U2-Pad2_ Net-_U5-Pad2_ Net-_X5-Pad4_ Net-_X10-Pad2_ 4_and
X5 Net-_U1-Pad10_ Net-_U2-Pad2_ Net-_U3-Pad2_ Net-_X5-Pad4_ Net-_X10-Pad1_ 4_and
X4 Net-_X1-Pad1_ Net-_U4-Pad2_ Net-_U5-Pad2_ Net-_U1-Pad3_ Net-_X4-Pad5_ 4_and
X10 Net-_X10-Pad1_ Net-_X10-Pad2_ Net-_X10-Pad3_ Net-_X10-Pad4_ Net-_U1-Pad9_ 4_OR
X8 Net-_U1-Pad13_ Net-_U4-Pad2_ Net-_U5-Pad2_ Net-_X5-Pad4_ Net-_X10-Pad4_ 4_and
X7 Net-_U1-Pad12_ Net-_U4-Pad2_ Net-_U3-Pad2_ Net-_X5-Pad4_ Net-_X10-Pad3_ 4_and
U7 Net-_U1-Pad1_ Net-_X1-Pad1_ d_inverter
.end
