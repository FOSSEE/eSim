* C:\FOSSEE\eSim\library\SubcircuitLibrary\ca3080\ca3080.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/23/24 19:02:23

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
Q2  Net-_D2-Pad1_ Net-_D3-Pad2_ Net-_D3-Pad1_ eSim_PNP		
Q1  Net-_D2-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
Q5  Net-_D4-Pad1_ Net-_Q5-Pad2_ Net-_Q1-Pad3_ eSim_NPN		
Q6  Net-_Q11-Pad2_ Net-_D2-Pad2_ Net-_D3-Pad2_ eSim_PNP		
Q4  Net-_Q11-Pad2_ Net-_D2-Pad1_ Net-_D2-Pad2_ eSim_PNP		
D2  Net-_D2-Pad1_ Net-_D2-Pad2_ eSim_Diode		
D3  Net-_D3-Pad1_ Net-_D3-Pad2_ eSim_Diode		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q3  Net-_Q1-Pad3_ Net-_D1-Pad1_ Net-_D1-Pad2_ eSim_NPN		
Q8  Net-_Q10-Pad1_ Net-_D4-Pad1_ Net-_D4-Pad2_ eSim_PNP		
Q7  Net-_D4-Pad1_ Net-_D5-Pad2_ Net-_D3-Pad1_ eSim_PNP		
D4  Net-_D4-Pad1_ Net-_D4-Pad2_ eSim_Diode		
Q10  Net-_Q10-Pad1_ Net-_D4-Pad2_ Net-_D5-Pad2_ eSim_PNP		
D5  Net-_D3-Pad1_ Net-_D5-Pad2_ eSim_Diode		
D6  Net-_D6-Pad1_ Net-_D1-Pad2_ eSim_Diode		
Q9  Net-_Q11-Pad2_ Net-_D6-Pad1_ Net-_D1-Pad2_ eSim_NPN		
Q11  Net-_Q10-Pad1_ Net-_Q11-Pad2_ Net-_D6-Pad1_ eSim_NPN		
U1  ? Net-_Q1-Pad2_ Net-_Q5-Pad2_ Net-_D1-Pad2_ Net-_D1-Pad1_ Net-_Q10-Pad1_ Net-_D3-Pad1_ ? PORT		

.end
