* /home/vsduser/Downloads/eSim-2.3/library/SubcircuitLibrary/TG_D_Latch/TG_D_Latch.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Jun 23 11:13:51 2025

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
SC1  /D Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad4_ sky130_fd_pr__pfet_01v8		
SC2  /D /clk Net-_SC1-Pad3_ Net-_SC2-Pad4_ sky130_fd_pr__nfet_01v8		
SC4  Net-_SC3-Pad1_ Net-_SC1-Pad2_ Net-_SC1-Pad3_ Net-_SC1-Pad4_ sky130_fd_pr__pfet_01v8		
U1  /D /clk Net-_SC2-Pad4_ Net-_SC1-Pad4_ Net-_U1-Pad5_ Net-_SC1-Pad3_ PORT		
scmode1  SKY130mode		
SC3  Net-_SC3-Pad1_ /clk Net-_SC1-Pad3_ Net-_SC2-Pad4_ sky130_fd_pr__nfet_01v8		
X1  /clk Net-_SC1-Pad4_ Net-_SC2-Pad4_ Net-_SC1-Pad2_ CMOS_INVTR		
X2  Net-_SC1-Pad3_ Net-_SC1-Pad4_ Net-_SC2-Pad4_ Net-_U1-Pad5_ CMOS_INVTR		
X3  Net-_U1-Pad5_ Net-_SC1-Pad4_ Net-_SC2-Pad4_ Net-_SC3-Pad1_ CMOS_INVTR		

.end
