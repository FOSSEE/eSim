* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Jun  4 14:46:46 2015

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
R3  5 6 4.7k		
R4  7 0 1k		
R1  1 3 10k		
C1  8 1 0.01u		
R2  0 8 1Meg		
C2  0 8 5p		
C3  8 7 4p		
C4  8 6 2p		
C5  6 7 0.5p		
C6  7 0 2u		
C7  6 2 5u		
C8  2 0 6p		
R5  2 0 2.2k		
v2  5 0 dc		
*U1  3 vplot8_1		
*U2  2 vplot8_1		
v1  3 0 AC		
J1  6 8 7 NJF		

.end
